library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package DataPackage is
type t_data_array is array(natural range <>) of std_logic_vector(31 downto 0);
constant DATA : t_data_array(1760 - 1 downto 0) := (
    0 => X"00000000",
    1 => X"00000a89",
    2 => X"00000000",
    3 => X"00038a2f",
    4 => X"00000000",
    5 => X"00000a89",
    6 => X"000730c4",
    7 => X"000000fa",
    8 => X"00000000",
    9 => X"00000a89",
    10 => X"000760c9",
    11 => X"000000fa",
    12 => X"00000000",
    13 => X"00000a89",
    14 => X"0007a0cd",
    15 => X"000000fa",
    16 => X"00000000",
    17 => X"00000a89",
    18 => X"0007f0d2",
    19 => X"000000fa",
    20 => X"00000000",
    21 => X"00000a89",
    22 => X"000850d8",
    23 => X"000000fa",
    24 => X"00000000",
    25 => X"00000a89",
    26 => X"0008b0df",
    27 => X"000000fa",
    28 => X"00000000",
    29 => X"00000a89",
    30 => X"000930e7",
    31 => X"000000fa",
    32 => X"00000000",
    33 => X"00000a89",
    34 => X"0009c0f1",
    35 => X"000000fa",
    36 => X"00000000",
    37 => X"00000a89",
    38 => X"000a50fb",
    39 => X"000000fa",
    40 => X"00000000",
    41 => X"00000a89",
    42 => X"000af105",
    43 => X"000000fa",
    44 => X"00000000",
    45 => X"00000a89",
    46 => X"000b8110",
    47 => X"000000fa",
    48 => X"00000000",
    49 => X"00000a89",
    50 => X"000bf11a",
    51 => X"000000fa",
    52 => X"00000000",
    53 => X"00000a89",
    54 => X"000c5123",
    55 => X"000000fa",
    56 => X"00000000",
    57 => X"00000a89",
    58 => X"000c912b",
    59 => X"000000fa",
    60 => X"00000000",
    61 => X"00000a89",
    62 => X"000cd133",
    63 => X"000000fa",
    64 => X"00000000",
    65 => X"00000a89",
    66 => X"000d313f",
    67 => X"000000fa",
    68 => X"00000000",
    69 => X"00000a89",
    70 => X"000d914b",
    71 => X"000000fa",
    72 => X"00000000",
    73 => X"00000a89",
    74 => X"000e0158",
    75 => X"000000fa",
    76 => X"00000000",
    77 => X"00000a89",
    78 => X"000e8166",
    79 => X"000000fa",
    80 => X"00000000",
    81 => X"00000a89",
    82 => X"000f1173",
    83 => X"000000fa",
    84 => X"00000000",
    85 => X"00000a89",
    86 => X"000fa180",
    87 => X"000000fa",
    88 => X"00000000",
    89 => X"00000a89",
    90 => X"0010318e",
    91 => X"000000fa",
    92 => X"00000000",
    93 => X"00000a89",
    94 => X"0010c19c",
    95 => X"000000fa",
    96 => X"00000000",
    97 => X"00000a89",
    98 => X"001151ac",
    99 => X"000000fa",
    100 => X"00000000",
    101 => X"00000a89",
    102 => X"0011d1bc",
    103 => X"000000fa",
    104 => X"00000000",
    105 => X"00000a89",
    106 => X"001241cd",
    107 => X"000000fa",
    108 => X"00000000",
    109 => X"00000a89",
    110 => X"0012c1de",
    111 => X"000000fa",
    112 => X"00000000",
    113 => X"00000a89",
    114 => X"001341ef",
    115 => X"000000fa",
    116 => X"00000000",
    117 => X"00000a89",
    118 => X"0013e201",
    119 => X"000000fa",
    120 => X"00000000",
    121 => X"00000a89",
    122 => X"00149213",
    123 => X"000000fa",
    124 => X"00000000",
    125 => X"00000a89",
    126 => X"00154227",
    127 => X"000000fa",
    128 => X"00000000",
    129 => X"00000a89",
    130 => X"0015f23a",
    131 => X"000000fa",
    132 => X"00000000",
    133 => X"00000a89",
    134 => X"0016a24e",
    135 => X"000000fa",
    136 => X"00000000",
    137 => X"00000a89",
    138 => X"00175262",
    139 => X"000000fa",
    140 => X"00000000",
    141 => X"00000a89",
    142 => X"00180277",
    143 => X"000000fa",
    144 => X"00000000",
    145 => X"00000a89",
    146 => X"0018b28d",
    147 => X"000000fa",
    148 => X"00000000",
    149 => X"00000a89",
    150 => X"001962a2",
    151 => X"000000fa",
    152 => X"00000000",
    153 => X"00000a89",
    154 => X"001a22b8",
    155 => X"000000fa",
    156 => X"00000000",
    157 => X"00000a89",
    158 => X"001af2ce",
    159 => X"000000fa",
    160 => X"00000000",
    161 => X"00000a89",
    162 => X"001bc2e6",
    163 => X"000000fa",
    164 => X"00000000",
    165 => X"00000a89",
    166 => X"001c82fe",
    167 => X"000000fa",
    168 => X"00000000",
    169 => X"00000a89",
    170 => X"001d5316",
    171 => X"000000fa",
    172 => X"00000000",
    173 => X"00000a89",
    174 => X"001e232e",
    175 => X"000000fa",
    176 => X"00000000",
    177 => X"00000a89",
    178 => X"001ef347",
    179 => X"000000fa",
    180 => X"00000000",
    181 => X"00000a89",
    182 => X"001fc360",
    183 => X"000000fa",
    184 => X"00000000",
    185 => X"00000a89",
    186 => X"00209379",
    187 => X"000000fa",
    188 => X"00000000",
    189 => X"00000a89",
    190 => X"00216392",
    191 => X"000000fa",
    192 => X"00000000",
    193 => X"00000a89",
    194 => X"002243ac",
    195 => X"000000fa",
    196 => X"00000000",
    197 => X"00000a89",
    198 => X"002313c5",
    199 => X"000000fa",
    200 => X"00000000",
    201 => X"00000a89",
    202 => X"0023e3df",
    203 => X"000000fa",
    204 => X"00000000",
    205 => X"00000a89",
    206 => X"0024a3f9",
    207 => X"000000fa",
    208 => X"00000000",
    209 => X"00000a89",
    210 => X"00257414",
    211 => X"000000fa",
    212 => X"00000000",
    213 => X"00000a89",
    214 => X"0026442e",
    215 => X"000000fa",
    216 => X"00000000",
    217 => X"00000a89",
    218 => X"00270448",
    219 => X"000000fa",
    220 => X"00000000",
    221 => X"00000a89",
    222 => X"0027c462",
    223 => X"000000fa",
    224 => X"00000000",
    225 => X"00000a89",
    226 => X"0028847c",
    227 => X"000000fa",
    228 => X"00000000",
    229 => X"00000a89",
    230 => X"00293495",
    231 => X"000000fa",
    232 => X"00000000",
    233 => X"00000a89",
    234 => X"0029e4ae",
    235 => X"000000fa",
    236 => X"00000000",
    237 => X"00000a89",
    238 => X"002a94c7",
    239 => X"000000fa",
    240 => X"00000000",
    241 => X"00000a89",
    242 => X"002b34df",
    243 => X"000000fa",
    244 => X"00000000",
    245 => X"00000a89",
    246 => X"002bd4f6",
    247 => X"000000fa",
    248 => X"00000000",
    249 => X"00000a89",
    250 => X"002c650d",
    251 => X"000000fa",
    252 => X"00000000",
    253 => X"00000a89",
    254 => X"002cf522",
    255 => X"000000fa",
    256 => X"00000000",
    257 => X"00000a89",
    258 => X"002d7536",
    259 => X"000000fa",
    260 => X"00000000",
    261 => X"00000a89",
    262 => X"002de549",
    263 => X"000000fa",
    264 => X"00000000",
    265 => X"00000a89",
    266 => X"002e555a",
    267 => X"000000fa",
    268 => X"00000000",
    269 => X"00000a89",
    270 => X"002eb569",
    271 => X"000000fa",
    272 => X"00000000",
    273 => X"00000a89",
    274 => X"002f0576",
    275 => X"000000fa",
    276 => X"00000000",
    277 => X"00000a89",
    278 => X"002f4582",
    279 => X"000000fa",
    280 => X"00000000",
    281 => X"00000a89",
    282 => X"002f758a",
    283 => X"000000fa",
    284 => X"00000000",
    285 => X"00000a89",
    286 => X"002f9591",
    287 => X"000000fa",
    288 => X"00000000",
    289 => X"00000a89",
    290 => X"002fb595",
    291 => X"000000fa",
    292 => X"00000000",
    293 => X"00000a89",
    294 => X"002fb596",
    295 => X"000000fa",
    296 => X"00000000",
    297 => X"00000a89",
    298 => X"002fb595",
    299 => X"000000fa",
    300 => X"00000000",
    301 => X"00000a89",
    302 => X"002fa592",
    303 => X"000000fa",
    304 => X"00000000",
    305 => X"00000a89",
    306 => X"002f758b",
    307 => X"000000fa",
    308 => X"00000000",
    309 => X"00000a89",
    310 => X"002f4583",
    311 => X"000000fa",
    312 => X"00000000",
    313 => X"00000a89",
    314 => X"002f0578",
    315 => X"000000fa",
    316 => X"00000000",
    317 => X"00000a89",
    318 => X"002eb56b",
    319 => X"000000fa",
    320 => X"00000000",
    321 => X"00000a89",
    322 => X"002e655c",
    323 => X"000000fa",
    324 => X"00000000",
    325 => X"00000a89",
    326 => X"002df54b",
    327 => X"000000fa",
    328 => X"00000000",
    329 => X"00000a89",
    330 => X"002d8539",
    331 => X"000000fa",
    332 => X"00000000",
    333 => X"00000a89",
    334 => X"002d0525",
    335 => X"000000fa",
    336 => X"00000000",
    337 => X"00000a89",
    338 => X"002c7510",
    339 => X"000000fa",
    340 => X"00000000",
    341 => X"00000a89",
    342 => X"002be4f9",
    343 => X"000000fa",
    344 => X"00000000",
    345 => X"00000a89",
    346 => X"002b44e2",
    347 => X"000000fa",
    348 => X"00000000",
    349 => X"00000a89",
    350 => X"002aa4ca",
    351 => X"000000fa",
    352 => X"00000000",
    353 => X"00000a89",
    354 => X"002a04b2",
    355 => X"000000fa",
    356 => X"00000000",
    357 => X"00000a89",
    358 => X"00295499",
    359 => X"000000fa",
    360 => X"00000000",
    361 => X"00000a89",
    362 => X"0028a47f",
    363 => X"000000fa",
    364 => X"00000000",
    365 => X"00000a89",
    366 => X"0027e466",
    367 => X"000000fa",
    368 => X"00000000",
    369 => X"00000a89",
    370 => X"0027244c",
    371 => X"000000fa",
    372 => X"00000000",
    373 => X"00000a89",
    374 => X"00265432",
    375 => X"000000fa",
    376 => X"00000000",
    377 => X"00000a89",
    378 => X"00259417",
    379 => X"000000fa",
    380 => X"00000000",
    381 => X"00000a89",
    382 => X"0024c3fd",
    383 => X"000000fa",
    384 => X"00000000",
    385 => X"00000a89",
    386 => X"0023f3e3",
    387 => X"000000fa",
    388 => X"00000000",
    389 => X"00000a89",
    390 => X"002323c9",
    391 => X"000000fa",
    392 => X"00000000",
    393 => X"00000a89",
    394 => X"002253af",
    395 => X"000000fa",
    396 => X"00000000",
    397 => X"00000a89",
    398 => X"00218395",
    399 => X"000000fa",
    400 => X"00000000",
    401 => X"00000a89",
    402 => X"0020b37c",
    403 => X"000000fa",
    404 => X"00000000",
    405 => X"00000a89",
    406 => X"001fe363",
    407 => X"000000fa",
    408 => X"00000000",
    409 => X"00000a89",
    410 => X"001f134a",
    411 => X"000000fa",
    412 => X"00000000",
    413 => X"00000a89",
    414 => X"001e4332",
    415 => X"000000fa",
    416 => X"00000000",
    417 => X"00000a89",
    418 => X"001d7319",
    419 => X"000000fa",
    420 => X"00000000",
    421 => X"00000a89",
    422 => X"001ca301",
    423 => X"000000fa",
    424 => X"00000000",
    425 => X"00000a89",
    426 => X"001bd2e9",
    427 => X"000000fa",
    428 => X"00000000",
    429 => X"00000a89",
    430 => X"001b12d2",
    431 => X"000000fa",
    432 => X"00000000",
    433 => X"00000a89",
    434 => X"001a42bb",
    435 => X"000000fa",
    436 => X"00000000",
    437 => X"00000a89",
    438 => X"001982a5",
    439 => X"000000fa",
    440 => X"00000000",
    441 => X"00000a89",
    442 => X"0018c28f",
    443 => X"000000fa",
    444 => X"00000000",
    445 => X"00000a89",
    446 => X"0018127a",
    447 => X"000000fa",
    448 => X"00000000",
    449 => X"00000a89",
    450 => X"00176265",
    451 => X"000000fa",
    452 => X"00000000",
    453 => X"00000a89",
    454 => X"0016b251",
    455 => X"000000fa",
    456 => X"00000000",
    457 => X"00000a89",
    458 => X"0016023d",
    459 => X"000000fa",
    460 => X"00000000",
    461 => X"00000a89",
    462 => X"00155229",
    463 => X"000000fa",
    464 => X"00000000",
    465 => X"00000a89",
    466 => X"0014a216",
    467 => X"000000fa",
    468 => X"00000000",
    469 => X"00000a89",
    470 => X"00140203",
    471 => X"000000fa",
    472 => X"00000000",
    473 => X"00000a89",
    474 => X"001361f1",
    475 => X"000000fa",
    476 => X"00000000",
    477 => X"00000a89",
    478 => X"0012d1e0",
    479 => X"000000fa",
    480 => X"00000000",
    481 => X"00000a89",
    482 => X"001251cf",
    483 => X"000000fa",
    484 => X"00000000",
    485 => X"00000a89",
    486 => X"0011e1be",
    487 => X"000000fa",
    488 => X"00000000",
    489 => X"00000a89",
    490 => X"001161ae",
    491 => X"000000fa",
    492 => X"00000000",
    493 => X"00000a89",
    494 => X"0010d19e",
    495 => X"000000fa",
    496 => X"00000000",
    497 => X"00000a89",
    498 => X"00104190",
    499 => X"000000fa",
    500 => X"00000000",
    501 => X"00000a89",
    502 => X"000fb182",
    503 => X"000000fa",
    504 => X"00000000",
    505 => X"00000a89",
    506 => X"000f2175",
    507 => X"000000fa",
    508 => X"00000000",
    509 => X"00000a89",
    510 => X"000e9167",
    511 => X"000000fa",
    512 => X"00000000",
    513 => X"00000a89",
    514 => X"000e115a",
    515 => X"000000fa",
    516 => X"00000000",
    517 => X"00000a89",
    518 => X"000da14d",
    519 => X"000000fa",
    520 => X"00000000",
    521 => X"00000a89",
    522 => X"000d3140",
    523 => X"000000fa",
    524 => X"00000000",
    525 => X"00000a89",
    526 => X"000ce135",
    527 => X"000000fa",
    528 => X"00000000",
    529 => X"00000a89",
    530 => X"000c912c",
    531 => X"000000fa",
    532 => X"00000000",
    533 => X"00000a89",
    534 => X"000c6124",
    535 => X"000000fa",
    536 => X"00000000",
    537 => X"00000a89",
    538 => X"000c011b",
    539 => X"000000fa",
    540 => X"00000000",
    541 => X"00000a89",
    542 => X"000b9111",
    543 => X"000000fa",
    544 => X"00000000",
    545 => X"00000a89",
    546 => X"000b0107",
    547 => X"000000fa",
    548 => X"00000000",
    549 => X"00000a89",
    550 => X"000a60fc",
    551 => X"000000fa",
    552 => X"00000000",
    553 => X"00000a89",
    554 => X"0009d0f2",
    555 => X"000000fa",
    556 => X"00000000",
    557 => X"00000a89",
    558 => X"000940e9",
    559 => X"000000fa",
    560 => X"00000000",
    561 => X"00000a89",
    562 => X"0008c0e0",
    563 => X"000000fa",
    564 => X"00000000",
    565 => X"00000a89",
    566 => X"000860d9",
    567 => X"000000fa",
    568 => X"00000000",
    569 => X"00000a89",
    570 => X"000800d3",
    571 => X"000000fa",
    572 => X"00000000",
    573 => X"00000a89",
    574 => X"0007b0cd",
    575 => X"000000fa",
    576 => X"00000000",
    577 => X"00000a89",
    578 => X"000760ca",
    579 => X"000000fa",
    580 => X"00000000",
    581 => X"00000a89",
    582 => X"000730c5",
    583 => X"0001a209",
    584 => X"00000000",
    585 => X"00000a89",
    586 => X"00000000",
    587 => X"00704237",
    588 => X"00000000",
    589 => X"0000cffb",
    590 => X"00000000",
    591 => X"000000fa",
    592 => X"00000000",
    593 => X"0000cffb",
    594 => X"00000000",
    595 => X"000000fa",
    596 => X"00000000",
    597 => X"0000cffb",
    598 => X"00000000",
    599 => X"000000fa",
    600 => X"00000000",
    601 => X"0000cffb",
    602 => X"00000000",
    603 => X"000000fa",
    604 => X"00000000",
    605 => X"0000cffb",
    606 => X"00000000",
    607 => X"000000fa",
    608 => X"00000000",
    609 => X"0000cffb",
    610 => X"00000000",
    611 => X"000000fa",
    612 => X"00000000",
    613 => X"0000cffb",
    614 => X"00000000",
    615 => X"000000fa",
    616 => X"00000000",
    617 => X"0000cffb",
    618 => X"00000000",
    619 => X"000000fa",
    620 => X"00000000",
    621 => X"0000cffb",
    622 => X"00000000",
    623 => X"000000fa",
    624 => X"00000000",
    625 => X"0000cffb",
    626 => X"00000000",
    627 => X"000000fa",
    628 => X"00000000",
    629 => X"0000cffb",
    630 => X"00000000",
    631 => X"000000fa",
    632 => X"00000000",
    633 => X"0000cffb",
    634 => X"00000000",
    635 => X"000000fa",
    636 => X"00000000",
    637 => X"0000cffb",
    638 => X"00000000",
    639 => X"000000fa",
    640 => X"00000000",
    641 => X"0000cffb",
    642 => X"00000000",
    643 => X"000000fa",
    644 => X"00000000",
    645 => X"0000cffb",
    646 => X"00000000",
    647 => X"000000fa",
    648 => X"00000000",
    649 => X"0000cffb",
    650 => X"00000000",
    651 => X"000000fa",
    652 => X"00000000",
    653 => X"0000cffb",
    654 => X"00000000",
    655 => X"000000fa",
    656 => X"00000000",
    657 => X"0000cffb",
    658 => X"00000000",
    659 => X"000000fa",
    660 => X"00000000",
    661 => X"0000cffb",
    662 => X"00000000",
    663 => X"000000fa",
    664 => X"00000000",
    665 => X"0000cffb",
    666 => X"00000000",
    667 => X"000000fa",
    668 => X"00000000",
    669 => X"0000cffb",
    670 => X"00000000",
    671 => X"000000fa",
    672 => X"00000000",
    673 => X"0000cffb",
    674 => X"00000000",
    675 => X"000000fa",
    676 => X"00000000",
    677 => X"0000cffb",
    678 => X"00000000",
    679 => X"000000fa",
    680 => X"00000000",
    681 => X"0000cffb",
    682 => X"00000000",
    683 => X"000000fa",
    684 => X"00000000",
    685 => X"0000cffb",
    686 => X"00000000",
    687 => X"000000fa",
    688 => X"00000000",
    689 => X"0000cffb",
    690 => X"00000000",
    691 => X"000000fa",
    692 => X"00000000",
    693 => X"0000cffb",
    694 => X"00000000",
    695 => X"000000fa",
    696 => X"00000000",
    697 => X"0000cffb",
    698 => X"00000000",
    699 => X"000000fa",
    700 => X"00000000",
    701 => X"0000cffb",
    702 => X"00000000",
    703 => X"000000fa",
    704 => X"00000000",
    705 => X"0000cffb",
    706 => X"00000000",
    707 => X"000000fa",
    708 => X"00000000",
    709 => X"0000cffb",
    710 => X"00000000",
    711 => X"000000fa",
    712 => X"00000000",
    713 => X"0000cffb",
    714 => X"00000000",
    715 => X"000000fa",
    716 => X"00000000",
    717 => X"0000cffb",
    718 => X"00000000",
    719 => X"000000fa",
    720 => X"00000000",
    721 => X"0000cffb",
    722 => X"00000000",
    723 => X"000000fa",
    724 => X"00000000",
    725 => X"0000cffb",
    726 => X"00000000",
    727 => X"000000fa",
    728 => X"00000000",
    729 => X"0000cffb",
    730 => X"00000000",
    731 => X"000000fa",
    732 => X"00000000",
    733 => X"0000cffb",
    734 => X"00000000",
    735 => X"000000fa",
    736 => X"00000000",
    737 => X"0000cffb",
    738 => X"00000000",
    739 => X"000000fa",
    740 => X"00000000",
    741 => X"0000cffb",
    742 => X"00000000",
    743 => X"000000fa",
    744 => X"00000000",
    745 => X"0000cffb",
    746 => X"00000000",
    747 => X"000000fa",
    748 => X"00000000",
    749 => X"0000cffb",
    750 => X"00000000",
    751 => X"000000fa",
    752 => X"00000000",
    753 => X"0000cffb",
    754 => X"00000000",
    755 => X"000000fa",
    756 => X"00000000",
    757 => X"0000cffb",
    758 => X"00000000",
    759 => X"000000fa",
    760 => X"00000000",
    761 => X"0000cffb",
    762 => X"00000000",
    763 => X"000000fa",
    764 => X"00000000",
    765 => X"0000cffb",
    766 => X"00000000",
    767 => X"000000fa",
    768 => X"00000000",
    769 => X"0000cffb",
    770 => X"00000000",
    771 => X"000000fa",
    772 => X"00000000",
    773 => X"0000cffb",
    774 => X"00000000",
    775 => X"000000fa",
    776 => X"00000000",
    777 => X"0000cffb",
    778 => X"00000000",
    779 => X"000000fa",
    780 => X"00000000",
    781 => X"0000cffb",
    782 => X"00000000",
    783 => X"000000fa",
    784 => X"00000000",
    785 => X"0000cffb",
    786 => X"00000000",
    787 => X"000000fa",
    788 => X"00000000",
    789 => X"0000cffb",
    790 => X"00000000",
    791 => X"000000fa",
    792 => X"00000000",
    793 => X"0000cffb",
    794 => X"00000000",
    795 => X"000000fa",
    796 => X"00000000",
    797 => X"0000cffb",
    798 => X"00000000",
    799 => X"000000fa",
    800 => X"00000000",
    801 => X"0000cffb",
    802 => X"00000000",
    803 => X"000000fa",
    804 => X"00000000",
    805 => X"0000cffb",
    806 => X"00000000",
    807 => X"000000fa",
    808 => X"00000000",
    809 => X"0000cffb",
    810 => X"00000000",
    811 => X"000000fa",
    812 => X"00000000",
    813 => X"0000cffb",
    814 => X"00000000",
    815 => X"000000fa",
    816 => X"00000000",
    817 => X"0000cffb",
    818 => X"00000000",
    819 => X"000000fa",
    820 => X"00000000",
    821 => X"0000cffb",
    822 => X"00000000",
    823 => X"000000fa",
    824 => X"00000000",
    825 => X"0000cffb",
    826 => X"00000000",
    827 => X"000000fa",
    828 => X"00000000",
    829 => X"0000cffb",
    830 => X"00000000",
    831 => X"000000fa",
    832 => X"00000000",
    833 => X"0000cffb",
    834 => X"00000000",
    835 => X"000000fa",
    836 => X"00000000",
    837 => X"0000cffb",
    838 => X"00000000",
    839 => X"000000fa",
    840 => X"00000000",
    841 => X"0000cffb",
    842 => X"00000000",
    843 => X"000000fa",
    844 => X"00000000",
    845 => X"0000cffb",
    846 => X"00000000",
    847 => X"000000fa",
    848 => X"00000000",
    849 => X"0000cffb",
    850 => X"00000000",
    851 => X"000000fa",
    852 => X"00000000",
    853 => X"0000cffb",
    854 => X"00000000",
    855 => X"000000fa",
    856 => X"00000000",
    857 => X"0000cffb",
    858 => X"00000000",
    859 => X"000000fa",
    860 => X"00000000",
    861 => X"0000cffb",
    862 => X"00000000",
    863 => X"000000fa",
    864 => X"00000000",
    865 => X"0000cffb",
    866 => X"00000000",
    867 => X"000000fa",
    868 => X"00000000",
    869 => X"0000cffb",
    870 => X"00000000",
    871 => X"000000fa",
    872 => X"00000000",
    873 => X"0000cffb",
    874 => X"00000000",
    875 => X"000000fa",
    876 => X"00000000",
    877 => X"0000cffb",
    878 => X"00000000",
    879 => X"000000fa",
    880 => X"00000000",
    881 => X"0000cffb",
    882 => X"00000000",
    883 => X"000000fa",
    884 => X"00000000",
    885 => X"0000cffb",
    886 => X"00000000",
    887 => X"000000fa",
    888 => X"00000000",
    889 => X"0000cffb",
    890 => X"00000000",
    891 => X"000000fa",
    892 => X"00000000",
    893 => X"0000cffb",
    894 => X"00000000",
    895 => X"000000fa",
    896 => X"00000000",
    897 => X"0000cffb",
    898 => X"00000000",
    899 => X"000000fa",
    900 => X"00000000",
    901 => X"0000cffb",
    902 => X"00000000",
    903 => X"000000fa",
    904 => X"00000000",
    905 => X"0000cffb",
    906 => X"00000000",
    907 => X"000000fa",
    908 => X"00000000",
    909 => X"0000cffb",
    910 => X"00000000",
    911 => X"000000fa",
    912 => X"00000000",
    913 => X"0000cffb",
    914 => X"00000000",
    915 => X"000000fa",
    916 => X"00000000",
    917 => X"0000cffb",
    918 => X"00000000",
    919 => X"000000fa",
    920 => X"00000000",
    921 => X"0000cffb",
    922 => X"00000000",
    923 => X"000000fa",
    924 => X"00000000",
    925 => X"0000cffb",
    926 => X"00000000",
    927 => X"000000fa",
    928 => X"00000000",
    929 => X"0000cffb",
    930 => X"00000000",
    931 => X"000000fa",
    932 => X"00000000",
    933 => X"0000cffb",
    934 => X"00000000",
    935 => X"000000fa",
    936 => X"00000000",
    937 => X"0000cffb",
    938 => X"00000000",
    939 => X"000000fa",
    940 => X"00000000",
    941 => X"0000cffb",
    942 => X"00000000",
    943 => X"000000fa",
    944 => X"00000000",
    945 => X"0000cffb",
    946 => X"00000000",
    947 => X"000000fa",
    948 => X"00000000",
    949 => X"0000cffb",
    950 => X"00000000",
    951 => X"000000fa",
    952 => X"00000000",
    953 => X"0000cffb",
    954 => X"00000000",
    955 => X"000000fa",
    956 => X"00000000",
    957 => X"0000cffb",
    958 => X"00000000",
    959 => X"000000fa",
    960 => X"00000000",
    961 => X"0000cffb",
    962 => X"00000000",
    963 => X"000000fa",
    964 => X"00000000",
    965 => X"0000cffb",
    966 => X"00000000",
    967 => X"000000fa",
    968 => X"00000000",
    969 => X"0000cffb",
    970 => X"00000000",
    971 => X"000000fa",
    972 => X"00000000",
    973 => X"0000cffb",
    974 => X"00000000",
    975 => X"000000fa",
    976 => X"00000000",
    977 => X"0000cffb",
    978 => X"00000000",
    979 => X"000000fa",
    980 => X"00000000",
    981 => X"0000cffb",
    982 => X"00000000",
    983 => X"000000fa",
    984 => X"00000000",
    985 => X"0000cffb",
    986 => X"00000000",
    987 => X"000000fa",
    988 => X"00000000",
    989 => X"0000cffb",
    990 => X"00000000",
    991 => X"000000fa",
    992 => X"00000000",
    993 => X"0000cffb",
    994 => X"00000000",
    995 => X"000000fa",
    996 => X"00000000",
    997 => X"0000cffb",
    998 => X"00000000",
    999 => X"000000fa",
    1000 => X"00000000",
    1001 => X"0000cffb",
    1002 => X"00000000",
    1003 => X"000000fa",
    1004 => X"00000000",
    1005 => X"0000cffb",
    1006 => X"00000000",
    1007 => X"000000fa",
    1008 => X"00000000",
    1009 => X"0000cffb",
    1010 => X"00000000",
    1011 => X"000000fa",
    1012 => X"00000000",
    1013 => X"0000cffb",
    1014 => X"00000000",
    1015 => X"000000fa",
    1016 => X"00000000",
    1017 => X"0000cffb",
    1018 => X"00000000",
    1019 => X"000000fa",
    1020 => X"00000000",
    1021 => X"0000cffb",
    1022 => X"00000000",
    1023 => X"000000fa",
    1024 => X"00000000",
    1025 => X"0000cffb",
    1026 => X"00000000",
    1027 => X"000000fa",
    1028 => X"00000000",
    1029 => X"0000cffb",
    1030 => X"00000000",
    1031 => X"000000fa",
    1032 => X"00000000",
    1033 => X"0000cffb",
    1034 => X"00000000",
    1035 => X"000000fa",
    1036 => X"00000000",
    1037 => X"0000cffb",
    1038 => X"00000000",
    1039 => X"000000fa",
    1040 => X"00000000",
    1041 => X"0000cffb",
    1042 => X"00000000",
    1043 => X"000000fa",
    1044 => X"00000000",
    1045 => X"0000cffb",
    1046 => X"00000000",
    1047 => X"000000fa",
    1048 => X"00000000",
    1049 => X"0000cffb",
    1050 => X"00000000",
    1051 => X"000000fa",
    1052 => X"00000000",
    1053 => X"0000cffb",
    1054 => X"00000000",
    1055 => X"000000fa",
    1056 => X"00000000",
    1057 => X"0000cffb",
    1058 => X"00000000",
    1059 => X"000000fa",
    1060 => X"00000000",
    1061 => X"0000cffb",
    1062 => X"00000000",
    1063 => X"000000fa",
    1064 => X"00000000",
    1065 => X"0000cffb",
    1066 => X"00000000",
    1067 => X"000000fa",
    1068 => X"00000000",
    1069 => X"0000cffb",
    1070 => X"00000000",
    1071 => X"000000fa",
    1072 => X"00000000",
    1073 => X"0000cffb",
    1074 => X"00000000",
    1075 => X"000000fa",
    1076 => X"00000000",
    1077 => X"0000cffb",
    1078 => X"00000000",
    1079 => X"000000fa",
    1080 => X"00000000",
    1081 => X"0000cffb",
    1082 => X"00000000",
    1083 => X"000000fa",
    1084 => X"00000000",
    1085 => X"0000cffb",
    1086 => X"00000000",
    1087 => X"000000fa",
    1088 => X"00000000",
    1089 => X"0000cffb",
    1090 => X"00000000",
    1091 => X"000000fa",
    1092 => X"00000000",
    1093 => X"0000cffb",
    1094 => X"00000000",
    1095 => X"000000fa",
    1096 => X"00000000",
    1097 => X"0000cffb",
    1098 => X"00000000",
    1099 => X"000000fa",
    1100 => X"00000000",
    1101 => X"0000cffb",
    1102 => X"00000000",
    1103 => X"000000fa",
    1104 => X"00000000",
    1105 => X"0000cffb",
    1106 => X"00000000",
    1107 => X"000000fa",
    1108 => X"00000000",
    1109 => X"0000cffb",
    1110 => X"00000000",
    1111 => X"000000fa",
    1112 => X"00000000",
    1113 => X"0000cffb",
    1114 => X"00000000",
    1115 => X"000000fa",
    1116 => X"00000000",
    1117 => X"0000cffb",
    1118 => X"00000000",
    1119 => X"000000fa",
    1120 => X"00000000",
    1121 => X"0000cffb",
    1122 => X"00000000",
    1123 => X"000000fa",
    1124 => X"00000000",
    1125 => X"0000cffb",
    1126 => X"00000000",
    1127 => X"000000fa",
    1128 => X"00000000",
    1129 => X"0000cffb",
    1130 => X"00000000",
    1131 => X"000000fa",
    1132 => X"00000000",
    1133 => X"0000cffb",
    1134 => X"00000000",
    1135 => X"000000fa",
    1136 => X"00000000",
    1137 => X"0000cffb",
    1138 => X"00000000",
    1139 => X"000000fa",
    1140 => X"00000000",
    1141 => X"0000cffb",
    1142 => X"00000000",
    1143 => X"000000fa",
    1144 => X"00000000",
    1145 => X"0000cffb",
    1146 => X"00000000",
    1147 => X"000000fa",
    1148 => X"00000000",
    1149 => X"0000cffb",
    1150 => X"00000000",
    1151 => X"000000fa",
    1152 => X"00000000",
    1153 => X"0000cffb",
    1154 => X"00000000",
    1155 => X"000000fa",
    1156 => X"00000000",
    1157 => X"0000cffb",
    1158 => X"00000000",
    1159 => X"000000fa",
    1160 => X"00000000",
    1161 => X"0000cffb",
    1162 => X"00000000",
    1163 => X"000000fa",
    1164 => X"00000000",
    1165 => X"0000cffb",
    1166 => X"00000000",
    1167 => X"0001a209",
    1168 => X"00000000",
    1169 => X"0000cffb",
    1170 => X"00000000",
    1171 => X"00704237",
    1172 => X"00000000",
    1173 => X"0001956c",
    1174 => X"00000000",
    1175 => X"000000fa",
    1176 => X"00000000",
    1177 => X"0001956c",
    1178 => X"00000000",
    1179 => X"000000fa",
    1180 => X"00000000",
    1181 => X"0001956c",
    1182 => X"00000000",
    1183 => X"000000fa",
    1184 => X"00000000",
    1185 => X"0001956c",
    1186 => X"00000000",
    1187 => X"000000fa",
    1188 => X"00000000",
    1189 => X"0001956c",
    1190 => X"00000000",
    1191 => X"000000fa",
    1192 => X"00000000",
    1193 => X"0001956c",
    1194 => X"00000000",
    1195 => X"000000fa",
    1196 => X"00000000",
    1197 => X"0001956c",
    1198 => X"00000000",
    1199 => X"000000fa",
    1200 => X"00000000",
    1201 => X"0001956c",
    1202 => X"00000000",
    1203 => X"000000fa",
    1204 => X"00000000",
    1205 => X"0001956c",
    1206 => X"00000000",
    1207 => X"000000fa",
    1208 => X"00000000",
    1209 => X"0001956c",
    1210 => X"00000000",
    1211 => X"000000fa",
    1212 => X"00000000",
    1213 => X"0001956c",
    1214 => X"00000000",
    1215 => X"000000fa",
    1216 => X"00000000",
    1217 => X"0001956c",
    1218 => X"00000000",
    1219 => X"000000fa",
    1220 => X"00000000",
    1221 => X"0001956c",
    1222 => X"00000000",
    1223 => X"000000fa",
    1224 => X"00000000",
    1225 => X"0001956c",
    1226 => X"00000000",
    1227 => X"000000fa",
    1228 => X"00000000",
    1229 => X"0001956c",
    1230 => X"00000000",
    1231 => X"000000fa",
    1232 => X"00000000",
    1233 => X"0001956c",
    1234 => X"00000000",
    1235 => X"000000fa",
    1236 => X"00000000",
    1237 => X"0001956c",
    1238 => X"00000000",
    1239 => X"000000fa",
    1240 => X"00000000",
    1241 => X"0001956c",
    1242 => X"00000000",
    1243 => X"000000fa",
    1244 => X"00000000",
    1245 => X"0001956c",
    1246 => X"00000000",
    1247 => X"000000fa",
    1248 => X"00000000",
    1249 => X"0001956c",
    1250 => X"00000000",
    1251 => X"000000fa",
    1252 => X"00000000",
    1253 => X"0001956c",
    1254 => X"00000000",
    1255 => X"000000fa",
    1256 => X"00000000",
    1257 => X"0001956c",
    1258 => X"00000000",
    1259 => X"000000fa",
    1260 => X"00000000",
    1261 => X"0001956c",
    1262 => X"00000000",
    1263 => X"000000fa",
    1264 => X"00000000",
    1265 => X"0001956c",
    1266 => X"00000000",
    1267 => X"000000fa",
    1268 => X"00000000",
    1269 => X"0001956c",
    1270 => X"00000000",
    1271 => X"000000fa",
    1272 => X"00000000",
    1273 => X"0001956c",
    1274 => X"00000000",
    1275 => X"000000fa",
    1276 => X"00000000",
    1277 => X"0001956c",
    1278 => X"00000000",
    1279 => X"000000fa",
    1280 => X"00000000",
    1281 => X"0001956c",
    1282 => X"00000000",
    1283 => X"000000fa",
    1284 => X"00000000",
    1285 => X"0001956c",
    1286 => X"00000000",
    1287 => X"000000fa",
    1288 => X"00000000",
    1289 => X"0001956c",
    1290 => X"00000000",
    1291 => X"000000fa",
    1292 => X"00000000",
    1293 => X"0001956c",
    1294 => X"00000000",
    1295 => X"000000fa",
    1296 => X"00000000",
    1297 => X"0001956c",
    1298 => X"00000000",
    1299 => X"000000fa",
    1300 => X"00000000",
    1301 => X"0001956c",
    1302 => X"00000000",
    1303 => X"000000fa",
    1304 => X"00000000",
    1305 => X"0001956c",
    1306 => X"00000000",
    1307 => X"000000fa",
    1308 => X"00000000",
    1309 => X"0001956c",
    1310 => X"00000000",
    1311 => X"000000fa",
    1312 => X"00000000",
    1313 => X"0001956c",
    1314 => X"00000000",
    1315 => X"000000fa",
    1316 => X"00000000",
    1317 => X"0001956c",
    1318 => X"00000000",
    1319 => X"000000fa",
    1320 => X"00000000",
    1321 => X"0001956c",
    1322 => X"00000000",
    1323 => X"000000fa",
    1324 => X"00000000",
    1325 => X"0001956c",
    1326 => X"00000000",
    1327 => X"000000fa",
    1328 => X"00000000",
    1329 => X"0001956c",
    1330 => X"00000000",
    1331 => X"000000fa",
    1332 => X"00000000",
    1333 => X"0001956c",
    1334 => X"00000000",
    1335 => X"000000fa",
    1336 => X"00000000",
    1337 => X"0001956c",
    1338 => X"00000000",
    1339 => X"000000fa",
    1340 => X"00000000",
    1341 => X"0001956c",
    1342 => X"00000000",
    1343 => X"000000fa",
    1344 => X"00000000",
    1345 => X"0001956c",
    1346 => X"00000000",
    1347 => X"000000fa",
    1348 => X"00000000",
    1349 => X"0001956c",
    1350 => X"00000000",
    1351 => X"000000fa",
    1352 => X"00000000",
    1353 => X"0001956c",
    1354 => X"00000000",
    1355 => X"000000fa",
    1356 => X"00000000",
    1357 => X"0001956c",
    1358 => X"00000000",
    1359 => X"000000fa",
    1360 => X"00000000",
    1361 => X"0001956c",
    1362 => X"00000000",
    1363 => X"000000fa",
    1364 => X"00000000",
    1365 => X"0001956c",
    1366 => X"00000000",
    1367 => X"000000fa",
    1368 => X"00000000",
    1369 => X"0001956c",
    1370 => X"00000000",
    1371 => X"000000fa",
    1372 => X"00000000",
    1373 => X"0001956c",
    1374 => X"00000000",
    1375 => X"000000fa",
    1376 => X"00000000",
    1377 => X"0001956c",
    1378 => X"00000000",
    1379 => X"000000fa",
    1380 => X"00000000",
    1381 => X"0001956c",
    1382 => X"00000000",
    1383 => X"000000fa",
    1384 => X"00000000",
    1385 => X"0001956c",
    1386 => X"00000000",
    1387 => X"000000fa",
    1388 => X"00000000",
    1389 => X"0001956c",
    1390 => X"00000000",
    1391 => X"000000fa",
    1392 => X"00000000",
    1393 => X"0001956c",
    1394 => X"00000000",
    1395 => X"000000fa",
    1396 => X"00000000",
    1397 => X"0001956c",
    1398 => X"00000000",
    1399 => X"000000fa",
    1400 => X"00000000",
    1401 => X"0001956c",
    1402 => X"00000000",
    1403 => X"000000fa",
    1404 => X"00000000",
    1405 => X"0001956c",
    1406 => X"00000000",
    1407 => X"000000fa",
    1408 => X"00000000",
    1409 => X"0001956c",
    1410 => X"00000000",
    1411 => X"000000fa",
    1412 => X"00000000",
    1413 => X"0001956c",
    1414 => X"00000000",
    1415 => X"000000fa",
    1416 => X"00000000",
    1417 => X"0001956c",
    1418 => X"00000000",
    1419 => X"000000fa",
    1420 => X"00000000",
    1421 => X"0001956c",
    1422 => X"00000000",
    1423 => X"000000fa",
    1424 => X"00000000",
    1425 => X"0001956c",
    1426 => X"00000000",
    1427 => X"000000fa",
    1428 => X"00000000",
    1429 => X"0001956c",
    1430 => X"00000000",
    1431 => X"000000fa",
    1432 => X"00000000",
    1433 => X"0001956c",
    1434 => X"00000000",
    1435 => X"000000fa",
    1436 => X"00000000",
    1437 => X"0001956c",
    1438 => X"00000000",
    1439 => X"000000fa",
    1440 => X"00000000",
    1441 => X"0001956c",
    1442 => X"00000000",
    1443 => X"000000fa",
    1444 => X"00000000",
    1445 => X"0001956c",
    1446 => X"00000000",
    1447 => X"000000fa",
    1448 => X"00000000",
    1449 => X"0001956c",
    1450 => X"00000000",
    1451 => X"000000fa",
    1452 => X"00000000",
    1453 => X"0001956c",
    1454 => X"00000000",
    1455 => X"000000fa",
    1456 => X"00000000",
    1457 => X"0001956c",
    1458 => X"00000000",
    1459 => X"000000fa",
    1460 => X"00000000",
    1461 => X"0001956c",
    1462 => X"00000000",
    1463 => X"000000fa",
    1464 => X"00000000",
    1465 => X"0001956c",
    1466 => X"00000000",
    1467 => X"000000fa",
    1468 => X"00000000",
    1469 => X"0001956c",
    1470 => X"00000000",
    1471 => X"000000fa",
    1472 => X"00000000",
    1473 => X"0001956c",
    1474 => X"00000000",
    1475 => X"000000fa",
    1476 => X"00000000",
    1477 => X"0001956c",
    1478 => X"00000000",
    1479 => X"000000fa",
    1480 => X"00000000",
    1481 => X"0001956c",
    1482 => X"00000000",
    1483 => X"000000fa",
    1484 => X"00000000",
    1485 => X"0001956c",
    1486 => X"00000000",
    1487 => X"000000fa",
    1488 => X"00000000",
    1489 => X"0001956c",
    1490 => X"00000000",
    1491 => X"000000fa",
    1492 => X"00000000",
    1493 => X"0001956c",
    1494 => X"00000000",
    1495 => X"000000fa",
    1496 => X"00000000",
    1497 => X"0001956c",
    1498 => X"00000000",
    1499 => X"000000fa",
    1500 => X"00000000",
    1501 => X"0001956c",
    1502 => X"00000000",
    1503 => X"000000fa",
    1504 => X"00000000",
    1505 => X"0001956c",
    1506 => X"00000000",
    1507 => X"000000fa",
    1508 => X"00000000",
    1509 => X"0001956c",
    1510 => X"00000000",
    1511 => X"000000fa",
    1512 => X"00000000",
    1513 => X"0001956c",
    1514 => X"00000000",
    1515 => X"000000fa",
    1516 => X"00000000",
    1517 => X"0001956c",
    1518 => X"00000000",
    1519 => X"000000fa",
    1520 => X"00000000",
    1521 => X"0001956c",
    1522 => X"00000000",
    1523 => X"000000fa",
    1524 => X"00000000",
    1525 => X"0001956c",
    1526 => X"00000000",
    1527 => X"000000fa",
    1528 => X"00000000",
    1529 => X"0001956c",
    1530 => X"00000000",
    1531 => X"000000fa",
    1532 => X"00000000",
    1533 => X"0001956c",
    1534 => X"00000000",
    1535 => X"000000fa",
    1536 => X"00000000",
    1537 => X"0001956c",
    1538 => X"00000000",
    1539 => X"000000fa",
    1540 => X"00000000",
    1541 => X"0001956c",
    1542 => X"00000000",
    1543 => X"000000fa",
    1544 => X"00000000",
    1545 => X"0001956c",
    1546 => X"00000000",
    1547 => X"000000fa",
    1548 => X"00000000",
    1549 => X"0001956c",
    1550 => X"00000000",
    1551 => X"000000fa",
    1552 => X"00000000",
    1553 => X"0001956c",
    1554 => X"00000000",
    1555 => X"000000fa",
    1556 => X"00000000",
    1557 => X"0001956c",
    1558 => X"00000000",
    1559 => X"000000fa",
    1560 => X"00000000",
    1561 => X"0001956c",
    1562 => X"00000000",
    1563 => X"000000fa",
    1564 => X"00000000",
    1565 => X"0001956c",
    1566 => X"00000000",
    1567 => X"000000fa",
    1568 => X"00000000",
    1569 => X"0001956c",
    1570 => X"00000000",
    1571 => X"000000fa",
    1572 => X"00000000",
    1573 => X"0001956c",
    1574 => X"00000000",
    1575 => X"000000fa",
    1576 => X"00000000",
    1577 => X"0001956c",
    1578 => X"00000000",
    1579 => X"000000fa",
    1580 => X"00000000",
    1581 => X"0001956c",
    1582 => X"00000000",
    1583 => X"000000fa",
    1584 => X"00000000",
    1585 => X"0001956c",
    1586 => X"00000000",
    1587 => X"000000fa",
    1588 => X"00000000",
    1589 => X"0001956c",
    1590 => X"00000000",
    1591 => X"000000fa",
    1592 => X"00000000",
    1593 => X"0001956c",
    1594 => X"00000000",
    1595 => X"000000fa",
    1596 => X"00000000",
    1597 => X"0001956c",
    1598 => X"00000000",
    1599 => X"000000fa",
    1600 => X"00000000",
    1601 => X"0001956c",
    1602 => X"00000000",
    1603 => X"000000fa",
    1604 => X"00000000",
    1605 => X"0001956c",
    1606 => X"00000000",
    1607 => X"000000fa",
    1608 => X"00000000",
    1609 => X"0001956c",
    1610 => X"00000000",
    1611 => X"000000fa",
    1612 => X"00000000",
    1613 => X"0001956c",
    1614 => X"00000000",
    1615 => X"000000fa",
    1616 => X"00000000",
    1617 => X"0001956c",
    1618 => X"00000000",
    1619 => X"000000fa",
    1620 => X"00000000",
    1621 => X"0001956c",
    1622 => X"00000000",
    1623 => X"000000fa",
    1624 => X"00000000",
    1625 => X"0001956c",
    1626 => X"00000000",
    1627 => X"000000fa",
    1628 => X"00000000",
    1629 => X"0001956c",
    1630 => X"00000000",
    1631 => X"000000fa",
    1632 => X"00000000",
    1633 => X"0001956c",
    1634 => X"00000000",
    1635 => X"000000fa",
    1636 => X"00000000",
    1637 => X"0001956c",
    1638 => X"00000000",
    1639 => X"000000fa",
    1640 => X"00000000",
    1641 => X"0001956c",
    1642 => X"00000000",
    1643 => X"000000fa",
    1644 => X"00000000",
    1645 => X"0001956c",
    1646 => X"00000000",
    1647 => X"000000fa",
    1648 => X"00000000",
    1649 => X"0001956c",
    1650 => X"00000000",
    1651 => X"000000fa",
    1652 => X"00000000",
    1653 => X"0001956c",
    1654 => X"00000000",
    1655 => X"000000fa",
    1656 => X"00000000",
    1657 => X"0001956c",
    1658 => X"00000000",
    1659 => X"000000fa",
    1660 => X"00000000",
    1661 => X"0001956c",
    1662 => X"00000000",
    1663 => X"000000fa",
    1664 => X"00000000",
    1665 => X"0001956c",
    1666 => X"00000000",
    1667 => X"000000fa",
    1668 => X"00000000",
    1669 => X"0001956c",
    1670 => X"00000000",
    1671 => X"000000fa",
    1672 => X"00000000",
    1673 => X"0001956c",
    1674 => X"00000000",
    1675 => X"000000fa",
    1676 => X"00000000",
    1677 => X"0001956c",
    1678 => X"00000000",
    1679 => X"000000fa",
    1680 => X"00000000",
    1681 => X"0001956c",
    1682 => X"00000000",
    1683 => X"000000fa",
    1684 => X"00000000",
    1685 => X"0001956c",
    1686 => X"00000000",
    1687 => X"000000fa",
    1688 => X"00000000",
    1689 => X"0001956c",
    1690 => X"00000000",
    1691 => X"000000fa",
    1692 => X"00000000",
    1693 => X"0001956c",
    1694 => X"00000000",
    1695 => X"000000fa",
    1696 => X"00000000",
    1697 => X"0001956c",
    1698 => X"00000000",
    1699 => X"000000fa",
    1700 => X"00000000",
    1701 => X"0001956c",
    1702 => X"00000000",
    1703 => X"000000fa",
    1704 => X"00000000",
    1705 => X"0001956c",
    1706 => X"00000000",
    1707 => X"000000fa",
    1708 => X"00000000",
    1709 => X"0001956c",
    1710 => X"00000000",
    1711 => X"000000fa",
    1712 => X"00000000",
    1713 => X"0001956c",
    1714 => X"00000000",
    1715 => X"000000fa",
    1716 => X"00000000",
    1717 => X"0001956c",
    1718 => X"00000000",
    1719 => X"000000fa",
    1720 => X"00000000",
    1721 => X"0001956c",
    1722 => X"00000000",
    1723 => X"000000fa",
    1724 => X"00000000",
    1725 => X"0001956c",
    1726 => X"00000000",
    1727 => X"000000fa",
    1728 => X"00000000",
    1729 => X"0001956c",
    1730 => X"00000000",
    1731 => X"000000fa",
    1732 => X"00000000",
    1733 => X"0001956c",
    1734 => X"00000000",
    1735 => X"000000fa",
    1736 => X"00000000",
    1737 => X"0001956c",
    1738 => X"00000000",
    1739 => X"000000fa",
    1740 => X"00000000",
    1741 => X"0001956c",
    1742 => X"00000000",
    1743 => X"000000fa",
    1744 => X"00000000",
    1745 => X"0001956c",
    1746 => X"00000000",
    1747 => X"000000fa",
    1748 => X"00000000",
    1749 => X"0001956c",
    1750 => X"00000000",
    1751 => X"0001a209",
    1752 => X"00000000",
    1753 => X"0001956c",
    1754 => X"00000000",
    1755 => X"000003e8",
    1756 => X"00000000",
    1757 => X"0001956c",
    1758 => X"00000000",
    1759 => X"00000000");
end DataPackage;
