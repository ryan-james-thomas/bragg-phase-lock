library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package DataPackage is
type t_data_array is array(natural range <>) of std_logic_vector(31 downto 0);
constant DATA : t_data_array(4008 - 1 downto 0) := (
    0 => X"00000000",
    1 => X"0000d1b7",
    2 => X"00000000",
    3 => X"000000fa",
    4 => X"00000000",
    5 => X"0000d1b7",
    6 => X"00000000",
    7 => X"000000fa",
    8 => X"00000000",
    9 => X"0000d1b7",
    10 => X"00000000",
    11 => X"000000fa",
    12 => X"00000000",
    13 => X"0000d1b7",
    14 => X"00000000",
    15 => X"000000fa",
    16 => X"00000000",
    17 => X"0000d1b7",
    18 => X"00000001",
    19 => X"000000fa",
    20 => X"00000000",
    21 => X"0000d1b7",
    22 => X"00000001",
    23 => X"000000fa",
    24 => X"00000000",
    25 => X"0000d1b7",
    26 => X"00000001",
    27 => X"000000fa",
    28 => X"00000000",
    29 => X"0000d1b7",
    30 => X"00000002",
    31 => X"000000fa",
    32 => X"00000000",
    33 => X"0000d1b7",
    34 => X"00000002",
    35 => X"000000fa",
    36 => X"00000000",
    37 => X"0000d1b7",
    38 => X"00000003",
    39 => X"000000fa",
    40 => X"00000000",
    41 => X"0000d1b7",
    42 => X"00000004",
    43 => X"000000fa",
    44 => X"00000000",
    45 => X"0000d1b7",
    46 => X"00000004",
    47 => X"000000fa",
    48 => X"00000000",
    49 => X"0000d1b7",
    50 => X"00000005",
    51 => X"000000fa",
    52 => X"00000000",
    53 => X"0000d1b7",
    54 => X"00000006",
    55 => X"000000fa",
    56 => X"00000000",
    57 => X"0000d1b7",
    58 => X"00000007",
    59 => X"000000fa",
    60 => X"00000000",
    61 => X"0000d1b7",
    62 => X"00000008",
    63 => X"000000fa",
    64 => X"00000000",
    65 => X"0000d1b7",
    66 => X"00000009",
    67 => X"000000fa",
    68 => X"00000000",
    69 => X"0000d1b7",
    70 => X"0000000b",
    71 => X"000000fa",
    72 => X"00000000",
    73 => X"0000d1b7",
    74 => X"0000000c",
    75 => X"000000fa",
    76 => X"00000000",
    77 => X"0000d1b7",
    78 => X"0000000d",
    79 => X"000000fa",
    80 => X"00000000",
    81 => X"0000d1b7",
    82 => X"0000000f",
    83 => X"000000fa",
    84 => X"00000000",
    85 => X"0000d1b7",
    86 => X"00000010",
    87 => X"000000fa",
    88 => X"00000000",
    89 => X"0000d1b7",
    90 => X"00000012",
    91 => X"000000fa",
    92 => X"00000000",
    93 => X"0000d1b7",
    94 => X"00000013",
    95 => X"000000fa",
    96 => X"00000000",
    97 => X"0000d1b7",
    98 => X"00000015",
    99 => X"000000fa",
    100 => X"00000000",
    101 => X"0000d1b7",
    102 => X"00000017",
    103 => X"000000fa",
    104 => X"00000000",
    105 => X"0000d1b7",
    106 => X"00000019",
    107 => X"000000fa",
    108 => X"00000000",
    109 => X"0000d1b7",
    110 => X"0000001a",
    111 => X"000000fa",
    112 => X"00000000",
    113 => X"0000d1b7",
    114 => X"0000001c",
    115 => X"000000fa",
    116 => X"00000000",
    117 => X"0000d1b7",
    118 => X"0000001f",
    119 => X"000000fa",
    120 => X"00000000",
    121 => X"0000d1b7",
    122 => X"00000021",
    123 => X"000000fa",
    124 => X"00000000",
    125 => X"0000d1b7",
    126 => X"00000023",
    127 => X"000000fa",
    128 => X"00000000",
    129 => X"0000d1b7",
    130 => X"00000025",
    131 => X"000000fa",
    132 => X"00000000",
    133 => X"0000d1b7",
    134 => X"00000027",
    135 => X"000000fa",
    136 => X"00000000",
    137 => X"0000d1b7",
    138 => X"0000002a",
    139 => X"000000fa",
    140 => X"00000000",
    141 => X"0000d1b7",
    142 => X"0000002c",
    143 => X"000000fa",
    144 => X"00000000",
    145 => X"0000d1b7",
    146 => X"0000002f",
    147 => X"000000fa",
    148 => X"00000000",
    149 => X"0000d1b7",
    150 => X"00000032",
    151 => X"000000fa",
    152 => X"00000000",
    153 => X"0000d1b7",
    154 => X"00000034",
    155 => X"000000fa",
    156 => X"00000000",
    157 => X"0000d1b7",
    158 => X"00000037",
    159 => X"000000fa",
    160 => X"00000000",
    161 => X"0000d1b7",
    162 => X"0000003a",
    163 => X"000000fa",
    164 => X"00000000",
    165 => X"0000d1b7",
    166 => X"0000003d",
    167 => X"000000fa",
    168 => X"00000000",
    169 => X"0000d1b7",
    170 => X"00000040",
    171 => X"000000fa",
    172 => X"00000000",
    173 => X"0000d1b7",
    174 => X"00000043",
    175 => X"000000fa",
    176 => X"00000000",
    177 => X"0000d1b7",
    178 => X"00000046",
    179 => X"000000fa",
    180 => X"00000000",
    181 => X"0000d1b7",
    182 => X"00000049",
    183 => X"000000fa",
    184 => X"00000000",
    185 => X"0000d1b7",
    186 => X"0000004c",
    187 => X"000000fa",
    188 => X"00000000",
    189 => X"0000d1b7",
    190 => X"00000050",
    191 => X"000000fa",
    192 => X"00000000",
    193 => X"0000d1b7",
    194 => X"00000053",
    195 => X"000000fa",
    196 => X"00000000",
    197 => X"0000d1b7",
    198 => X"00000057",
    199 => X"000000fa",
    200 => X"00000000",
    201 => X"0000d1b7",
    202 => X"0000005a",
    203 => X"000000fa",
    204 => X"00000000",
    205 => X"0000d1b7",
    206 => X"0000005e",
    207 => X"000000fa",
    208 => X"00000000",
    209 => X"0000d1b7",
    210 => X"00000061",
    211 => X"000000fa",
    212 => X"00000000",
    213 => X"0000d1b7",
    214 => X"00000065",
    215 => X"000000fa",
    216 => X"00000000",
    217 => X"0000d1b7",
    218 => X"00000069",
    219 => X"000000fa",
    220 => X"00000000",
    221 => X"0000d1b7",
    222 => X"0000006d",
    223 => X"000000fa",
    224 => X"00000000",
    225 => X"0000d1b7",
    226 => X"00000071",
    227 => X"000000fa",
    228 => X"00000000",
    229 => X"0000d1b7",
    230 => X"00000075",
    231 => X"000000fa",
    232 => X"00000000",
    233 => X"0000d1b7",
    234 => X"00000079",
    235 => X"000000fa",
    236 => X"00000000",
    237 => X"0000d1b7",
    238 => X"0000007d",
    239 => X"000000fa",
    240 => X"00000000",
    241 => X"0000d1b7",
    242 => X"00000081",
    243 => X"000000fa",
    244 => X"00000000",
    245 => X"0000d1b7",
    246 => X"00000086",
    247 => X"000000fa",
    248 => X"00000000",
    249 => X"0000d1b7",
    250 => X"0000008a",
    251 => X"000000fa",
    252 => X"00000000",
    253 => X"0000d1b7",
    254 => X"0000008e",
    255 => X"000000fa",
    256 => X"00000000",
    257 => X"0000d1b7",
    258 => X"00000093",
    259 => X"000000fa",
    260 => X"00000000",
    261 => X"0000d1b7",
    262 => X"00000098",
    263 => X"000000fa",
    264 => X"00000000",
    265 => X"0000d1b7",
    266 => X"0000009c",
    267 => X"000000fa",
    268 => X"00000000",
    269 => X"0000d1b7",
    270 => X"000000a1",
    271 => X"000000fa",
    272 => X"00000000",
    273 => X"0000d1b7",
    274 => X"000000a6",
    275 => X"000000fa",
    276 => X"00000000",
    277 => X"0000d1b7",
    278 => X"000000aa",
    279 => X"000000fa",
    280 => X"00000000",
    281 => X"0000d1b7",
    282 => X"000000af",
    283 => X"000000fa",
    284 => X"00000000",
    285 => X"0000d1b7",
    286 => X"000000b4",
    287 => X"000000fa",
    288 => X"00000000",
    289 => X"0000d1b7",
    290 => X"000000b9",
    291 => X"000000fa",
    292 => X"00000000",
    293 => X"0000d1b7",
    294 => X"000000be",
    295 => X"000000fa",
    296 => X"00000000",
    297 => X"0000d1b7",
    298 => X"000000c4",
    299 => X"000000fa",
    300 => X"00000000",
    301 => X"0000d1b7",
    302 => X"000000c9",
    303 => X"000000fa",
    304 => X"00000000",
    305 => X"0000d1b7",
    306 => X"000000ce",
    307 => X"000000fa",
    308 => X"00000000",
    309 => X"0000d1b7",
    310 => X"000000d3",
    311 => X"000000fa",
    312 => X"00000000",
    313 => X"0000d1b7",
    314 => X"000000d9",
    315 => X"000000fa",
    316 => X"00000000",
    317 => X"0000d1b7",
    318 => X"000000de",
    319 => X"000000fa",
    320 => X"00000000",
    321 => X"0000d1b7",
    322 => X"000000e4",
    323 => X"000000fa",
    324 => X"00000000",
    325 => X"0000d1b7",
    326 => X"000000ea",
    327 => X"000000fa",
    328 => X"00000000",
    329 => X"0000d1b7",
    330 => X"000000ef",
    331 => X"000000fa",
    332 => X"00000000",
    333 => X"0000d1b7",
    334 => X"000000f5",
    335 => X"000000fa",
    336 => X"00000000",
    337 => X"0000d1b7",
    338 => X"000000fb",
    339 => X"000000fa",
    340 => X"00000000",
    341 => X"0000d1b7",
    342 => X"00000101",
    343 => X"000000fa",
    344 => X"00000000",
    345 => X"0000d1b7",
    346 => X"00000107",
    347 => X"000000fa",
    348 => X"00000000",
    349 => X"0000d1b7",
    350 => X"0000010d",
    351 => X"000000fa",
    352 => X"00000000",
    353 => X"0000d1b7",
    354 => X"00000113",
    355 => X"000000fa",
    356 => X"00000000",
    357 => X"0000d1b7",
    358 => X"00000119",
    359 => X"000000fa",
    360 => X"00000000",
    361 => X"0000d1b7",
    362 => X"0000011f",
    363 => X"000000fa",
    364 => X"00000000",
    365 => X"0000d1b7",
    366 => X"00000125",
    367 => X"000000fa",
    368 => X"00000000",
    369 => X"0000d1b7",
    370 => X"0000012b",
    371 => X"000000fa",
    372 => X"00000000",
    373 => X"0000d1b7",
    374 => X"00000132",
    375 => X"000000fa",
    376 => X"00000000",
    377 => X"0000d1b7",
    378 => X"00000138",
    379 => X"000000fa",
    380 => X"00000000",
    381 => X"0000d1b7",
    382 => X"0000013f",
    383 => X"000000fa",
    384 => X"00000000",
    385 => X"0000d1b7",
    386 => X"00000145",
    387 => X"000000fa",
    388 => X"00000000",
    389 => X"0000d1b7",
    390 => X"0000014c",
    391 => X"000000fa",
    392 => X"00000000",
    393 => X"0000d1b7",
    394 => X"00000152",
    395 => X"000000fa",
    396 => X"00000000",
    397 => X"0000d1b7",
    398 => X"00000159",
    399 => X"000000fa",
    400 => X"00000000",
    401 => X"0000d1b7",
    402 => X"00000160",
    403 => X"000000fa",
    404 => X"00000000",
    405 => X"0000d1b7",
    406 => X"00000167",
    407 => X"000000fa",
    408 => X"00000000",
    409 => X"0000d1b7",
    410 => X"0000016e",
    411 => X"000000fa",
    412 => X"00000000",
    413 => X"0000d1b7",
    414 => X"00000175",
    415 => X"000000fa",
    416 => X"00000000",
    417 => X"0000d1b7",
    418 => X"0000017c",
    419 => X"000000fa",
    420 => X"00000000",
    421 => X"0000d1b7",
    422 => X"00000183",
    423 => X"000000fa",
    424 => X"00000000",
    425 => X"0000d1b7",
    426 => X"0000018a",
    427 => X"000000fa",
    428 => X"00000000",
    429 => X"0000d1b7",
    430 => X"00000191",
    431 => X"000000fa",
    432 => X"00000000",
    433 => X"0000d1b7",
    434 => X"00000198",
    435 => X"000000fa",
    436 => X"00000000",
    437 => X"0000d1b7",
    438 => X"000001a0",
    439 => X"000000fa",
    440 => X"00000000",
    441 => X"0000d1b7",
    442 => X"000001a7",
    443 => X"000000fa",
    444 => X"00000000",
    445 => X"0000d1b7",
    446 => X"000001ae",
    447 => X"000000fa",
    448 => X"00000000",
    449 => X"0000d1b7",
    450 => X"000001b6",
    451 => X"000000fa",
    452 => X"00000000",
    453 => X"0000d1b7",
    454 => X"000001bd",
    455 => X"000000fa",
    456 => X"00000000",
    457 => X"0000d1b7",
    458 => X"000001c5",
    459 => X"000000fa",
    460 => X"00000000",
    461 => X"0000d1b7",
    462 => X"000001cc",
    463 => X"000000fa",
    464 => X"00000000",
    465 => X"0000d1b7",
    466 => X"000001d4",
    467 => X"000000fa",
    468 => X"00000000",
    469 => X"0000d1b7",
    470 => X"000001dc",
    471 => X"000000fa",
    472 => X"00000000",
    473 => X"0000d1b7",
    474 => X"000001e4",
    475 => X"000000fa",
    476 => X"00000000",
    477 => X"0000d1b7",
    478 => X"000001ec",
    479 => X"000000fa",
    480 => X"00000000",
    481 => X"0000d1b7",
    482 => X"000001f3",
    483 => X"000000fa",
    484 => X"00000000",
    485 => X"0000d1b7",
    486 => X"000001fb",
    487 => X"000000fa",
    488 => X"00000000",
    489 => X"0000d1b7",
    490 => X"00000203",
    491 => X"000000fa",
    492 => X"00000000",
    493 => X"0000d1b7",
    494 => X"0000020b",
    495 => X"000000fa",
    496 => X"00000000",
    497 => X"0000d1b7",
    498 => X"00000214",
    499 => X"000000fa",
    500 => X"00000000",
    501 => X"0000d1b7",
    502 => X"0000021c",
    503 => X"000000fa",
    504 => X"00000000",
    505 => X"0000d1b7",
    506 => X"00000224",
    507 => X"000000fa",
    508 => X"00000000",
    509 => X"0000d1b7",
    510 => X"0000022c",
    511 => X"000000fa",
    512 => X"00000000",
    513 => X"0000d1b7",
    514 => X"00000235",
    515 => X"000000fa",
    516 => X"00000000",
    517 => X"0000d1b7",
    518 => X"0000023d",
    519 => X"000000fa",
    520 => X"00000000",
    521 => X"0000d1b7",
    522 => X"00000245",
    523 => X"000000fa",
    524 => X"00000000",
    525 => X"0000d1b7",
    526 => X"0000024e",
    527 => X"000000fa",
    528 => X"00000000",
    529 => X"0000d1b7",
    530 => X"00000256",
    531 => X"000000fa",
    532 => X"00000000",
    533 => X"0000d1b7",
    534 => X"0000025f",
    535 => X"000000fa",
    536 => X"00000000",
    537 => X"0000d1b7",
    538 => X"00000267",
    539 => X"000000fa",
    540 => X"00000000",
    541 => X"0000d1b7",
    542 => X"00000270",
    543 => X"000000fa",
    544 => X"00000000",
    545 => X"0000d1b7",
    546 => X"00000279",
    547 => X"000000fa",
    548 => X"00000000",
    549 => X"0000d1b7",
    550 => X"00000282",
    551 => X"000000fa",
    552 => X"00000000",
    553 => X"0000d1b7",
    554 => X"0000028a",
    555 => X"000000fa",
    556 => X"00000000",
    557 => X"0000d1b7",
    558 => X"00000293",
    559 => X"000000fa",
    560 => X"00000000",
    561 => X"0000d1b7",
    562 => X"0000029c",
    563 => X"000000fa",
    564 => X"00000000",
    565 => X"0000d1b7",
    566 => X"000002a5",
    567 => X"000000fa",
    568 => X"00000000",
    569 => X"0000d1b7",
    570 => X"000002ae",
    571 => X"000000fa",
    572 => X"00000000",
    573 => X"0000d1b7",
    574 => X"000002b7",
    575 => X"000000fa",
    576 => X"00000000",
    577 => X"0000d1b7",
    578 => X"000002c0",
    579 => X"000000fa",
    580 => X"00000000",
    581 => X"0000d1b7",
    582 => X"000002c9",
    583 => X"000000fa",
    584 => X"00000000",
    585 => X"0000d1b7",
    586 => X"000002d2",
    587 => X"000000fa",
    588 => X"00000000",
    589 => X"0000d1b7",
    590 => X"000002dc",
    591 => X"000000fa",
    592 => X"00000000",
    593 => X"0000d1b7",
    594 => X"000002e5",
    595 => X"000000fa",
    596 => X"00000000",
    597 => X"0000d1b7",
    598 => X"000002ee",
    599 => X"000000fa",
    600 => X"00000000",
    601 => X"0000d1b7",
    602 => X"000002f8",
    603 => X"000000fa",
    604 => X"00000000",
    605 => X"0000d1b7",
    606 => X"00000301",
    607 => X"000000fa",
    608 => X"00000000",
    609 => X"0000d1b7",
    610 => X"0000030a",
    611 => X"000000fa",
    612 => X"00000000",
    613 => X"0000d1b7",
    614 => X"00000314",
    615 => X"000000fa",
    616 => X"00000000",
    617 => X"0000d1b7",
    618 => X"0000031d",
    619 => X"000000fa",
    620 => X"00000000",
    621 => X"0000d1b7",
    622 => X"00000327",
    623 => X"000000fa",
    624 => X"00000000",
    625 => X"0000d1b7",
    626 => X"00000331",
    627 => X"000000fa",
    628 => X"00000000",
    629 => X"0000d1b7",
    630 => X"0000033a",
    631 => X"000000fa",
    632 => X"00000000",
    633 => X"0000d1b7",
    634 => X"00000344",
    635 => X"000000fa",
    636 => X"00000000",
    637 => X"0000d1b7",
    638 => X"0000034e",
    639 => X"000000fa",
    640 => X"00000000",
    641 => X"0000d1b7",
    642 => X"00000357",
    643 => X"000000fa",
    644 => X"00000000",
    645 => X"0000d1b7",
    646 => X"00000361",
    647 => X"000000fa",
    648 => X"00000000",
    649 => X"0000d1b7",
    650 => X"0000036b",
    651 => X"000000fa",
    652 => X"00000000",
    653 => X"0000d1b7",
    654 => X"00000375",
    655 => X"000000fa",
    656 => X"00000000",
    657 => X"0000d1b7",
    658 => X"0000037f",
    659 => X"000000fa",
    660 => X"00000000",
    661 => X"0000d1b7",
    662 => X"00000389",
    663 => X"000000fa",
    664 => X"00000000",
    665 => X"0000d1b7",
    666 => X"00000393",
    667 => X"000000fa",
    668 => X"00000000",
    669 => X"0000d1b7",
    670 => X"0000039d",
    671 => X"000000fa",
    672 => X"00000000",
    673 => X"0000d1b7",
    674 => X"000003a7",
    675 => X"000000fa",
    676 => X"00000000",
    677 => X"0000d1b7",
    678 => X"000003b1",
    679 => X"000000fa",
    680 => X"00000000",
    681 => X"0000d1b7",
    682 => X"000003bb",
    683 => X"000000fa",
    684 => X"00000000",
    685 => X"0000d1b7",
    686 => X"000003c5",
    687 => X"000000fa",
    688 => X"00000000",
    689 => X"0000d1b7",
    690 => X"000003cf",
    691 => X"000000fa",
    692 => X"00000000",
    693 => X"0000d1b7",
    694 => X"000003da",
    695 => X"000000fa",
    696 => X"00000000",
    697 => X"0000d1b7",
    698 => X"000003e4",
    699 => X"000000fa",
    700 => X"00000000",
    701 => X"0000d1b7",
    702 => X"000003ee",
    703 => X"000000fa",
    704 => X"00000000",
    705 => X"0000d1b7",
    706 => X"000003f8",
    707 => X"000000fa",
    708 => X"00000000",
    709 => X"0000d1b7",
    710 => X"00000403",
    711 => X"000000fa",
    712 => X"00000000",
    713 => X"0000d1b7",
    714 => X"0000040d",
    715 => X"000000fa",
    716 => X"00000000",
    717 => X"0000d1b7",
    718 => X"00000418",
    719 => X"000000fa",
    720 => X"00000000",
    721 => X"0000d1b7",
    722 => X"00000422",
    723 => X"000000fa",
    724 => X"00000000",
    725 => X"0000d1b7",
    726 => X"0000042d",
    727 => X"000000fa",
    728 => X"00000000",
    729 => X"0000d1b7",
    730 => X"00000437",
    731 => X"000000fa",
    732 => X"00000000",
    733 => X"0000d1b7",
    734 => X"00000442",
    735 => X"000000fa",
    736 => X"00000000",
    737 => X"0000d1b7",
    738 => X"0000044c",
    739 => X"000000fa",
    740 => X"00000000",
    741 => X"0000d1b7",
    742 => X"00000457",
    743 => X"000000fa",
    744 => X"00000000",
    745 => X"0000d1b7",
    746 => X"00000462",
    747 => X"000000fa",
    748 => X"00000000",
    749 => X"0000d1b7",
    750 => X"0000046c",
    751 => X"000000fa",
    752 => X"00000000",
    753 => X"0000d1b7",
    754 => X"00000477",
    755 => X"000000fa",
    756 => X"00000000",
    757 => X"0000d1b7",
    758 => X"00000482",
    759 => X"000000fa",
    760 => X"00000000",
    761 => X"0000d1b7",
    762 => X"0000048c",
    763 => X"000000fa",
    764 => X"00000000",
    765 => X"0000d1b7",
    766 => X"00000497",
    767 => X"000000fa",
    768 => X"00000000",
    769 => X"0000d1b7",
    770 => X"000004a2",
    771 => X"000000fa",
    772 => X"00000000",
    773 => X"0000d1b7",
    774 => X"000004ad",
    775 => X"000000fa",
    776 => X"00000000",
    777 => X"0000d1b7",
    778 => X"000004b8",
    779 => X"000000fa",
    780 => X"00000000",
    781 => X"0000d1b7",
    782 => X"000004c3",
    783 => X"000000fa",
    784 => X"00000000",
    785 => X"0000d1b7",
    786 => X"000004cd",
    787 => X"000000fa",
    788 => X"00000000",
    789 => X"0000d1b7",
    790 => X"000004d8",
    791 => X"000000fa",
    792 => X"00000000",
    793 => X"0000d1b7",
    794 => X"000004e3",
    795 => X"000000fa",
    796 => X"00000000",
    797 => X"0000d1b7",
    798 => X"000004ee",
    799 => X"000000fa",
    800 => X"00000000",
    801 => X"0000d1b7",
    802 => X"000004f9",
    803 => X"000000fa",
    804 => X"00000000",
    805 => X"0000d1b7",
    806 => X"00000504",
    807 => X"000000fa",
    808 => X"00000000",
    809 => X"0000d1b7",
    810 => X"0000050f",
    811 => X"000000fa",
    812 => X"00000000",
    813 => X"0000d1b7",
    814 => X"0000051a",
    815 => X"000000fa",
    816 => X"00000000",
    817 => X"0000d1b7",
    818 => X"00000526",
    819 => X"000000fa",
    820 => X"00000000",
    821 => X"0000d1b7",
    822 => X"00000531",
    823 => X"000000fa",
    824 => X"00000000",
    825 => X"0000d1b7",
    826 => X"0000053c",
    827 => X"000000fa",
    828 => X"00000000",
    829 => X"0000d1b7",
    830 => X"00000547",
    831 => X"000000fa",
    832 => X"00000000",
    833 => X"0000d1b7",
    834 => X"00000552",
    835 => X"000000fa",
    836 => X"00000000",
    837 => X"0000d1b7",
    838 => X"0000055d",
    839 => X"000000fa",
    840 => X"00000000",
    841 => X"0000d1b7",
    842 => X"00000568",
    843 => X"000000fa",
    844 => X"00000000",
    845 => X"0000d1b7",
    846 => X"00000574",
    847 => X"000000fa",
    848 => X"00000000",
    849 => X"0000d1b7",
    850 => X"0000057f",
    851 => X"000000fa",
    852 => X"00000000",
    853 => X"0000d1b7",
    854 => X"0000058a",
    855 => X"000000fa",
    856 => X"00000000",
    857 => X"0000d1b7",
    858 => X"00000595",
    859 => X"000000fa",
    860 => X"00000000",
    861 => X"0000d1b7",
    862 => X"000005a1",
    863 => X"000000fa",
    864 => X"00000000",
    865 => X"0000d1b7",
    866 => X"000005ac",
    867 => X"000000fa",
    868 => X"00000000",
    869 => X"0000d1b7",
    870 => X"000005b7",
    871 => X"000000fa",
    872 => X"00000000",
    873 => X"0000d1b7",
    874 => X"000005c3",
    875 => X"000000fa",
    876 => X"00000000",
    877 => X"0000d1b7",
    878 => X"000005ce",
    879 => X"000000fa",
    880 => X"00000000",
    881 => X"0000d1b7",
    882 => X"000005d9",
    883 => X"000000fa",
    884 => X"00000000",
    885 => X"0000d1b7",
    886 => X"000005e5",
    887 => X"000000fa",
    888 => X"00000000",
    889 => X"0000d1b7",
    890 => X"000005f0",
    891 => X"000000fa",
    892 => X"00000000",
    893 => X"0000d1b7",
    894 => X"000005fc",
    895 => X"000000fa",
    896 => X"00000000",
    897 => X"0000d1b7",
    898 => X"00000607",
    899 => X"000000fa",
    900 => X"00000000",
    901 => X"0000d1b7",
    902 => X"00000612",
    903 => X"000000fa",
    904 => X"00000000",
    905 => X"0000d1b7",
    906 => X"0000061e",
    907 => X"000000fa",
    908 => X"00000000",
    909 => X"0000d1b7",
    910 => X"00000629",
    911 => X"000000fa",
    912 => X"00000000",
    913 => X"0000d1b7",
    914 => X"00000635",
    915 => X"000000fa",
    916 => X"00000000",
    917 => X"0000d1b7",
    918 => X"00000640",
    919 => X"000000fa",
    920 => X"00000000",
    921 => X"0000d1b7",
    922 => X"0000064c",
    923 => X"000000fa",
    924 => X"00000000",
    925 => X"0000d1b7",
    926 => X"00000657",
    927 => X"000000fa",
    928 => X"00000000",
    929 => X"0000d1b7",
    930 => X"00000663",
    931 => X"000000fa",
    932 => X"00000000",
    933 => X"0000d1b7",
    934 => X"0000066e",
    935 => X"000000fa",
    936 => X"00000000",
    937 => X"0000d1b7",
    938 => X"0000067a",
    939 => X"000000fa",
    940 => X"00000000",
    941 => X"0000d1b7",
    942 => X"00000685",
    943 => X"000000fa",
    944 => X"00000000",
    945 => X"0000d1b7",
    946 => X"00000691",
    947 => X"000000fa",
    948 => X"00000000",
    949 => X"0000d1b7",
    950 => X"0000069c",
    951 => X"000000fa",
    952 => X"00000000",
    953 => X"0000d1b7",
    954 => X"000006a8",
    955 => X"000000fa",
    956 => X"00000000",
    957 => X"0000d1b7",
    958 => X"000006b3",
    959 => X"000000fa",
    960 => X"00000000",
    961 => X"0000d1b7",
    962 => X"000006bf",
    963 => X"000000fa",
    964 => X"00000000",
    965 => X"0000d1b7",
    966 => X"000006cb",
    967 => X"000000fa",
    968 => X"00000000",
    969 => X"0000d1b7",
    970 => X"000006d6",
    971 => X"000000fa",
    972 => X"00000000",
    973 => X"0000d1b7",
    974 => X"000006e2",
    975 => X"000000fa",
    976 => X"00000000",
    977 => X"0000d1b7",
    978 => X"000006ed",
    979 => X"000000fa",
    980 => X"00000000",
    981 => X"0000d1b7",
    982 => X"000006f9",
    983 => X"000000fa",
    984 => X"00000000",
    985 => X"0000d1b7",
    986 => X"00000704",
    987 => X"000000fa",
    988 => X"00000000",
    989 => X"0000d1b7",
    990 => X"00000710",
    991 => X"000000fa",
    992 => X"00000000",
    993 => X"0000d1b7",
    994 => X"0000071c",
    995 => X"000000fa",
    996 => X"00000000",
    997 => X"0000d1b7",
    998 => X"00000727",
    999 => X"000000fa",
    1000 => X"00000000",
    1001 => X"0000d1b7",
    1002 => X"00000733",
    1003 => X"000000fa",
    1004 => X"00000000",
    1005 => X"0000d1b7",
    1006 => X"0000073e",
    1007 => X"000000fa",
    1008 => X"00000000",
    1009 => X"0000d1b7",
    1010 => X"0000074a",
    1011 => X"000000fa",
    1012 => X"00000000",
    1013 => X"0000d1b7",
    1014 => X"00000755",
    1015 => X"000000fa",
    1016 => X"00000000",
    1017 => X"0000d1b7",
    1018 => X"00000761",
    1019 => X"000000fa",
    1020 => X"00000000",
    1021 => X"0000d1b7",
    1022 => X"0000076d",
    1023 => X"000000fa",
    1024 => X"00000000",
    1025 => X"0000d1b7",
    1026 => X"00000778",
    1027 => X"000000fa",
    1028 => X"00000000",
    1029 => X"0000d1b7",
    1030 => X"00000784",
    1031 => X"000000fa",
    1032 => X"00000000",
    1033 => X"0000d1b7",
    1034 => X"0000078f",
    1035 => X"000000fa",
    1036 => X"00000000",
    1037 => X"0000d1b7",
    1038 => X"0000079b",
    1039 => X"000000fa",
    1040 => X"00000000",
    1041 => X"0000d1b7",
    1042 => X"000007a6",
    1043 => X"000000fa",
    1044 => X"00000000",
    1045 => X"0000d1b7",
    1046 => X"000007b2",
    1047 => X"000000fa",
    1048 => X"00000000",
    1049 => X"0000d1b7",
    1050 => X"000007be",
    1051 => X"000000fa",
    1052 => X"00000000",
    1053 => X"0000d1b7",
    1054 => X"000007c9",
    1055 => X"000000fa",
    1056 => X"00000000",
    1057 => X"0000d1b7",
    1058 => X"000007d5",
    1059 => X"000000fa",
    1060 => X"00000000",
    1061 => X"0000d1b7",
    1062 => X"000007e0",
    1063 => X"000000fa",
    1064 => X"00000000",
    1065 => X"0000d1b7",
    1066 => X"000007ec",
    1067 => X"000000fa",
    1068 => X"00000000",
    1069 => X"0000d1b7",
    1070 => X"000007f7",
    1071 => X"000000fa",
    1072 => X"00000000",
    1073 => X"0000d1b7",
    1074 => X"00000803",
    1075 => X"000000fa",
    1076 => X"00000000",
    1077 => X"0000d1b7",
    1078 => X"0000080e",
    1079 => X"000000fa",
    1080 => X"00000000",
    1081 => X"0000d1b7",
    1082 => X"0000081a",
    1083 => X"000000fa",
    1084 => X"00000000",
    1085 => X"0000d1b7",
    1086 => X"00000825",
    1087 => X"000000fa",
    1088 => X"00000000",
    1089 => X"0000d1b7",
    1090 => X"00000831",
    1091 => X"000000fa",
    1092 => X"00000000",
    1093 => X"0000d1b7",
    1094 => X"0000083c",
    1095 => X"000000fa",
    1096 => X"00000000",
    1097 => X"0000d1b7",
    1098 => X"00000848",
    1099 => X"000000fa",
    1100 => X"00000000",
    1101 => X"0000d1b7",
    1102 => X"00000853",
    1103 => X"000000fa",
    1104 => X"00000000",
    1105 => X"0000d1b7",
    1106 => X"0000085e",
    1107 => X"000000fa",
    1108 => X"00000000",
    1109 => X"0000d1b7",
    1110 => X"0000086a",
    1111 => X"000000fa",
    1112 => X"00000000",
    1113 => X"0000d1b7",
    1114 => X"00000875",
    1115 => X"000000fa",
    1116 => X"00000000",
    1117 => X"0000d1b7",
    1118 => X"00000881",
    1119 => X"000000fa",
    1120 => X"00000000",
    1121 => X"0000d1b7",
    1122 => X"0000088c",
    1123 => X"000000fa",
    1124 => X"00000000",
    1125 => X"0000d1b7",
    1126 => X"00000897",
    1127 => X"000000fa",
    1128 => X"00000000",
    1129 => X"0000d1b7",
    1130 => X"000008a3",
    1131 => X"000000fa",
    1132 => X"00000000",
    1133 => X"0000d1b7",
    1134 => X"000008ae",
    1135 => X"000000fa",
    1136 => X"00000000",
    1137 => X"0000d1b7",
    1138 => X"000008b9",
    1139 => X"000000fa",
    1140 => X"00000000",
    1141 => X"0000d1b7",
    1142 => X"000008c5",
    1143 => X"000000fa",
    1144 => X"00000000",
    1145 => X"0000d1b7",
    1146 => X"000008d0",
    1147 => X"000000fa",
    1148 => X"00000000",
    1149 => X"0000d1b7",
    1150 => X"000008db",
    1151 => X"000000fa",
    1152 => X"00000000",
    1153 => X"0000d1b7",
    1154 => X"000008e7",
    1155 => X"000000fa",
    1156 => X"00000000",
    1157 => X"0000d1b7",
    1158 => X"000008f2",
    1159 => X"000000fa",
    1160 => X"00000000",
    1161 => X"0000d1b7",
    1162 => X"000008fd",
    1163 => X"000000fa",
    1164 => X"00000000",
    1165 => X"0000d1b7",
    1166 => X"00000908",
    1167 => X"000000fa",
    1168 => X"00000000",
    1169 => X"0000d1b7",
    1170 => X"00000913",
    1171 => X"000000fa",
    1172 => X"00000000",
    1173 => X"0000d1b7",
    1174 => X"0000091f",
    1175 => X"000000fa",
    1176 => X"00000000",
    1177 => X"0000d1b7",
    1178 => X"0000092a",
    1179 => X"000000fa",
    1180 => X"00000000",
    1181 => X"0000d1b7",
    1182 => X"00000935",
    1183 => X"000000fa",
    1184 => X"00000000",
    1185 => X"0000d1b7",
    1186 => X"00000940",
    1187 => X"000000fa",
    1188 => X"00000000",
    1189 => X"0000d1b7",
    1190 => X"0000094b",
    1191 => X"000000fa",
    1192 => X"00000000",
    1193 => X"0000d1b7",
    1194 => X"00000956",
    1195 => X"000000fa",
    1196 => X"00000000",
    1197 => X"0000d1b7",
    1198 => X"00000961",
    1199 => X"000000fa",
    1200 => X"00000000",
    1201 => X"0000d1b7",
    1202 => X"0000096c",
    1203 => X"000000fa",
    1204 => X"00000000",
    1205 => X"0000d1b7",
    1206 => X"00000977",
    1207 => X"000000fa",
    1208 => X"00000000",
    1209 => X"0000d1b7",
    1210 => X"00000982",
    1211 => X"000000fa",
    1212 => X"00000000",
    1213 => X"0000d1b7",
    1214 => X"0000098d",
    1215 => X"000000fa",
    1216 => X"00000000",
    1217 => X"0000d1b7",
    1218 => X"00000998",
    1219 => X"000000fa",
    1220 => X"00000000",
    1221 => X"0000d1b7",
    1222 => X"000009a3",
    1223 => X"000000fa",
    1224 => X"00000000",
    1225 => X"0000d1b7",
    1226 => X"000009ae",
    1227 => X"000000fa",
    1228 => X"00000000",
    1229 => X"0000d1b7",
    1230 => X"000009b9",
    1231 => X"000000fa",
    1232 => X"00000000",
    1233 => X"0000d1b7",
    1234 => X"000009c4",
    1235 => X"000000fa",
    1236 => X"00000000",
    1237 => X"0000d1b7",
    1238 => X"000009ce",
    1239 => X"000000fa",
    1240 => X"00000000",
    1241 => X"0000d1b7",
    1242 => X"000009d9",
    1243 => X"000000fa",
    1244 => X"00000000",
    1245 => X"0000d1b7",
    1246 => X"000009e4",
    1247 => X"000000fa",
    1248 => X"00000000",
    1249 => X"0000d1b7",
    1250 => X"000009ef",
    1251 => X"000000fa",
    1252 => X"00000000",
    1253 => X"0000d1b7",
    1254 => X"000009f9",
    1255 => X"000000fa",
    1256 => X"00000000",
    1257 => X"0000d1b7",
    1258 => X"00000a04",
    1259 => X"000000fa",
    1260 => X"00000000",
    1261 => X"0000d1b7",
    1262 => X"00000a0f",
    1263 => X"000000fa",
    1264 => X"00000000",
    1265 => X"0000d1b7",
    1266 => X"00000a19",
    1267 => X"000000fa",
    1268 => X"00000000",
    1269 => X"0000d1b7",
    1270 => X"00000a24",
    1271 => X"000000fa",
    1272 => X"00000000",
    1273 => X"0000d1b7",
    1274 => X"00000a2e",
    1275 => X"000000fa",
    1276 => X"00000000",
    1277 => X"0000d1b7",
    1278 => X"00000a39",
    1279 => X"000000fa",
    1280 => X"00000000",
    1281 => X"0000d1b7",
    1282 => X"00000a43",
    1283 => X"000000fa",
    1284 => X"00000000",
    1285 => X"0000d1b7",
    1286 => X"00000a4e",
    1287 => X"000000fa",
    1288 => X"00000000",
    1289 => X"0000d1b7",
    1290 => X"00000a58",
    1291 => X"000000fa",
    1292 => X"00000000",
    1293 => X"0000d1b7",
    1294 => X"00000a63",
    1295 => X"000000fa",
    1296 => X"00000000",
    1297 => X"0000d1b7",
    1298 => X"00000a6d",
    1299 => X"000000fa",
    1300 => X"00000000",
    1301 => X"0000d1b7",
    1302 => X"00000a77",
    1303 => X"000000fa",
    1304 => X"00000000",
    1305 => X"0000d1b7",
    1306 => X"00000a82",
    1307 => X"000000fa",
    1308 => X"00000000",
    1309 => X"0000d1b7",
    1310 => X"00000a8c",
    1311 => X"000000fa",
    1312 => X"00000000",
    1313 => X"0000d1b7",
    1314 => X"00000a96",
    1315 => X"000000fa",
    1316 => X"00000000",
    1317 => X"0000d1b7",
    1318 => X"00000aa0",
    1319 => X"000000fa",
    1320 => X"00000000",
    1321 => X"0000d1b7",
    1322 => X"00000aab",
    1323 => X"000000fa",
    1324 => X"00000000",
    1325 => X"0000d1b7",
    1326 => X"00000ab5",
    1327 => X"000000fa",
    1328 => X"00000000",
    1329 => X"0000d1b7",
    1330 => X"00000abf",
    1331 => X"000000fa",
    1332 => X"00000000",
    1333 => X"0000d1b7",
    1334 => X"00000ac9",
    1335 => X"000000fa",
    1336 => X"00000000",
    1337 => X"0000d1b7",
    1338 => X"00000ad3",
    1339 => X"000000fa",
    1340 => X"00000000",
    1341 => X"0000d1b7",
    1342 => X"00000add",
    1343 => X"000000fa",
    1344 => X"00000000",
    1345 => X"0000d1b7",
    1346 => X"00000ae7",
    1347 => X"000000fa",
    1348 => X"00000000",
    1349 => X"0000d1b7",
    1350 => X"00000af1",
    1351 => X"000000fa",
    1352 => X"00000000",
    1353 => X"0000d1b7",
    1354 => X"00000afb",
    1355 => X"000000fa",
    1356 => X"00000000",
    1357 => X"0000d1b7",
    1358 => X"00000b04",
    1359 => X"000000fa",
    1360 => X"00000000",
    1361 => X"0000d1b7",
    1362 => X"00000b0e",
    1363 => X"000000fa",
    1364 => X"00000000",
    1365 => X"0000d1b7",
    1366 => X"00000b18",
    1367 => X"000000fa",
    1368 => X"00000000",
    1369 => X"0000d1b7",
    1370 => X"00000b22",
    1371 => X"000000fa",
    1372 => X"00000000",
    1373 => X"0000d1b7",
    1374 => X"00000b2b",
    1375 => X"000000fa",
    1376 => X"00000000",
    1377 => X"0000d1b7",
    1378 => X"00000b35",
    1379 => X"000000fa",
    1380 => X"00000000",
    1381 => X"0000d1b7",
    1382 => X"00000b3f",
    1383 => X"000000fa",
    1384 => X"00000000",
    1385 => X"0000d1b7",
    1386 => X"00000b48",
    1387 => X"000000fa",
    1388 => X"00000000",
    1389 => X"0000d1b7",
    1390 => X"00000b52",
    1391 => X"000000fa",
    1392 => X"00000000",
    1393 => X"0000d1b7",
    1394 => X"00000b5b",
    1395 => X"000000fa",
    1396 => X"00000000",
    1397 => X"0000d1b7",
    1398 => X"00000b65",
    1399 => X"000000fa",
    1400 => X"00000000",
    1401 => X"0000d1b7",
    1402 => X"00000b6e",
    1403 => X"000000fa",
    1404 => X"00000000",
    1405 => X"0000d1b7",
    1406 => X"00000b77",
    1407 => X"000000fa",
    1408 => X"00000000",
    1409 => X"0000d1b7",
    1410 => X"00000b81",
    1411 => X"000000fa",
    1412 => X"00000000",
    1413 => X"0000d1b7",
    1414 => X"00000b8a",
    1415 => X"000000fa",
    1416 => X"00000000",
    1417 => X"0000d1b7",
    1418 => X"00000b93",
    1419 => X"000000fa",
    1420 => X"00000000",
    1421 => X"0000d1b7",
    1422 => X"00000b9c",
    1423 => X"000000fa",
    1424 => X"00000000",
    1425 => X"0000d1b7",
    1426 => X"00000ba5",
    1427 => X"000000fa",
    1428 => X"00000000",
    1429 => X"0000d1b7",
    1430 => X"00000bae",
    1431 => X"000000fa",
    1432 => X"00000000",
    1433 => X"0000d1b7",
    1434 => X"00000bb7",
    1435 => X"000000fa",
    1436 => X"00000000",
    1437 => X"0000d1b7",
    1438 => X"00000bc0",
    1439 => X"000000fa",
    1440 => X"00000000",
    1441 => X"0000d1b7",
    1442 => X"00000bc9",
    1443 => X"000000fa",
    1444 => X"00000000",
    1445 => X"0000d1b7",
    1446 => X"00000bd2",
    1447 => X"000000fa",
    1448 => X"00000000",
    1449 => X"0000d1b7",
    1450 => X"00000bdb",
    1451 => X"000000fa",
    1452 => X"00000000",
    1453 => X"0000d1b7",
    1454 => X"00000be4",
    1455 => X"000000fa",
    1456 => X"00000000",
    1457 => X"0000d1b7",
    1458 => X"00000bed",
    1459 => X"000000fa",
    1460 => X"00000000",
    1461 => X"0000d1b7",
    1462 => X"00000bf5",
    1463 => X"000000fa",
    1464 => X"00000000",
    1465 => X"0000d1b7",
    1466 => X"00000bfe",
    1467 => X"000000fa",
    1468 => X"00000000",
    1469 => X"0000d1b7",
    1470 => X"00000c07",
    1471 => X"000000fa",
    1472 => X"00000000",
    1473 => X"0000d1b7",
    1474 => X"00000c0f",
    1475 => X"000000fa",
    1476 => X"00000000",
    1477 => X"0000d1b7",
    1478 => X"00000c18",
    1479 => X"000000fa",
    1480 => X"00000000",
    1481 => X"0000d1b7",
    1482 => X"00000c20",
    1483 => X"000000fa",
    1484 => X"00000000",
    1485 => X"0000d1b7",
    1486 => X"00000c29",
    1487 => X"000000fa",
    1488 => X"00000000",
    1489 => X"0000d1b7",
    1490 => X"00000c31",
    1491 => X"000000fa",
    1492 => X"00000000",
    1493 => X"0000d1b7",
    1494 => X"00000c39",
    1495 => X"000000fa",
    1496 => X"00000000",
    1497 => X"0000d1b7",
    1498 => X"00000c42",
    1499 => X"000000fa",
    1500 => X"00000000",
    1501 => X"0000d1b7",
    1502 => X"00000c4a",
    1503 => X"000000fa",
    1504 => X"00000000",
    1505 => X"0000d1b7",
    1506 => X"00000c52",
    1507 => X"000000fa",
    1508 => X"00000000",
    1509 => X"0000d1b7",
    1510 => X"00000c5a",
    1511 => X"000000fa",
    1512 => X"00000000",
    1513 => X"0000d1b7",
    1514 => X"00000c62",
    1515 => X"000000fa",
    1516 => X"00000000",
    1517 => X"0000d1b7",
    1518 => X"00000c6a",
    1519 => X"000000fa",
    1520 => X"00000000",
    1521 => X"0000d1b7",
    1522 => X"00000c72",
    1523 => X"000000fa",
    1524 => X"00000000",
    1525 => X"0000d1b7",
    1526 => X"00000c7a",
    1527 => X"000000fa",
    1528 => X"00000000",
    1529 => X"0000d1b7",
    1530 => X"00000c82",
    1531 => X"000000fa",
    1532 => X"00000000",
    1533 => X"0000d1b7",
    1534 => X"00000c8a",
    1535 => X"000000fa",
    1536 => X"00000000",
    1537 => X"0000d1b7",
    1538 => X"00000c91",
    1539 => X"000000fa",
    1540 => X"00000000",
    1541 => X"0000d1b7",
    1542 => X"00000c99",
    1543 => X"000000fa",
    1544 => X"00000000",
    1545 => X"0000d1b7",
    1546 => X"00000ca1",
    1547 => X"000000fa",
    1548 => X"00000000",
    1549 => X"0000d1b7",
    1550 => X"00000ca8",
    1551 => X"000000fa",
    1552 => X"00000000",
    1553 => X"0000d1b7",
    1554 => X"00000cb0",
    1555 => X"000000fa",
    1556 => X"00000000",
    1557 => X"0000d1b7",
    1558 => X"00000cb7",
    1559 => X"000000fa",
    1560 => X"00000000",
    1561 => X"0000d1b7",
    1562 => X"00000cbf",
    1563 => X"000000fa",
    1564 => X"00000000",
    1565 => X"0000d1b7",
    1566 => X"00000cc6",
    1567 => X"000000fa",
    1568 => X"00000000",
    1569 => X"0000d1b7",
    1570 => X"00000ccd",
    1571 => X"000000fa",
    1572 => X"00000000",
    1573 => X"0000d1b7",
    1574 => X"00000cd5",
    1575 => X"000000fa",
    1576 => X"00000000",
    1577 => X"0000d1b7",
    1578 => X"00000cdc",
    1579 => X"000000fa",
    1580 => X"00000000",
    1581 => X"0000d1b7",
    1582 => X"00000ce3",
    1583 => X"000000fa",
    1584 => X"00000000",
    1585 => X"0000d1b7",
    1586 => X"00000cea",
    1587 => X"000000fa",
    1588 => X"00000000",
    1589 => X"0000d1b7",
    1590 => X"00000cf1",
    1591 => X"000000fa",
    1592 => X"00000000",
    1593 => X"0000d1b7",
    1594 => X"00000cf8",
    1595 => X"000000fa",
    1596 => X"00000000",
    1597 => X"0000d1b7",
    1598 => X"00000cff",
    1599 => X"000000fa",
    1600 => X"00000000",
    1601 => X"0000d1b7",
    1602 => X"00000d06",
    1603 => X"000000fa",
    1604 => X"00000000",
    1605 => X"0000d1b7",
    1606 => X"00000d0c",
    1607 => X"000000fa",
    1608 => X"00000000",
    1609 => X"0000d1b7",
    1610 => X"00000d13",
    1611 => X"000000fa",
    1612 => X"00000000",
    1613 => X"0000d1b7",
    1614 => X"00000d1a",
    1615 => X"000000fa",
    1616 => X"00000000",
    1617 => X"0000d1b7",
    1618 => X"00000d20",
    1619 => X"000000fa",
    1620 => X"00000000",
    1621 => X"0000d1b7",
    1622 => X"00000d27",
    1623 => X"000000fa",
    1624 => X"00000000",
    1625 => X"0000d1b7",
    1626 => X"00000d2d",
    1627 => X"000000fa",
    1628 => X"00000000",
    1629 => X"0000d1b7",
    1630 => X"00000d34",
    1631 => X"000000fa",
    1632 => X"00000000",
    1633 => X"0000d1b7",
    1634 => X"00000d3a",
    1635 => X"000000fa",
    1636 => X"00000000",
    1637 => X"0000d1b7",
    1638 => X"00000d40",
    1639 => X"000000fa",
    1640 => X"00000000",
    1641 => X"0000d1b7",
    1642 => X"00000d47",
    1643 => X"000000fa",
    1644 => X"00000000",
    1645 => X"0000d1b7",
    1646 => X"00000d4d",
    1647 => X"000000fa",
    1648 => X"00000000",
    1649 => X"0000d1b7",
    1650 => X"00000d53",
    1651 => X"000000fa",
    1652 => X"00000000",
    1653 => X"0000d1b7",
    1654 => X"00000d59",
    1655 => X"000000fa",
    1656 => X"00000000",
    1657 => X"0000d1b7",
    1658 => X"00000d5f",
    1659 => X"000000fa",
    1660 => X"00000000",
    1661 => X"0000d1b7",
    1662 => X"00000d65",
    1663 => X"000000fa",
    1664 => X"00000000",
    1665 => X"0000d1b7",
    1666 => X"00000d6b",
    1667 => X"000000fa",
    1668 => X"00000000",
    1669 => X"0000d1b7",
    1670 => X"00000d71",
    1671 => X"000000fa",
    1672 => X"00000000",
    1673 => X"0000d1b7",
    1674 => X"00000d76",
    1675 => X"000000fa",
    1676 => X"00000000",
    1677 => X"0000d1b7",
    1678 => X"00000d7c",
    1679 => X"000000fa",
    1680 => X"00000000",
    1681 => X"0000d1b7",
    1682 => X"00000d82",
    1683 => X"000000fa",
    1684 => X"00000000",
    1685 => X"0000d1b7",
    1686 => X"00000d87",
    1687 => X"000000fa",
    1688 => X"00000000",
    1689 => X"0000d1b7",
    1690 => X"00000d8d",
    1691 => X"000000fa",
    1692 => X"00000000",
    1693 => X"0000d1b7",
    1694 => X"00000d92",
    1695 => X"000000fa",
    1696 => X"00000000",
    1697 => X"0000d1b7",
    1698 => X"00000d97",
    1699 => X"000000fa",
    1700 => X"00000000",
    1701 => X"0000d1b7",
    1702 => X"00000d9d",
    1703 => X"000000fa",
    1704 => X"00000000",
    1705 => X"0000d1b7",
    1706 => X"00000da2",
    1707 => X"000000fa",
    1708 => X"00000000",
    1709 => X"0000d1b7",
    1710 => X"00000da7",
    1711 => X"000000fa",
    1712 => X"00000000",
    1713 => X"0000d1b7",
    1714 => X"00000dac",
    1715 => X"000000fa",
    1716 => X"00000000",
    1717 => X"0000d1b7",
    1718 => X"00000db1",
    1719 => X"000000fa",
    1720 => X"00000000",
    1721 => X"0000d1b7",
    1722 => X"00000db6",
    1723 => X"000000fa",
    1724 => X"00000000",
    1725 => X"0000d1b7",
    1726 => X"00000dbb",
    1727 => X"000000fa",
    1728 => X"00000000",
    1729 => X"0000d1b7",
    1730 => X"00000dc0",
    1731 => X"000000fa",
    1732 => X"00000000",
    1733 => X"0000d1b7",
    1734 => X"00000dc5",
    1735 => X"000000fa",
    1736 => X"00000000",
    1737 => X"0000d1b7",
    1738 => X"00000dc9",
    1739 => X"000000fa",
    1740 => X"00000000",
    1741 => X"0000d1b7",
    1742 => X"00000dce",
    1743 => X"000000fa",
    1744 => X"00000000",
    1745 => X"0000d1b7",
    1746 => X"00000dd3",
    1747 => X"000000fa",
    1748 => X"00000000",
    1749 => X"0000d1b7",
    1750 => X"00000dd7",
    1751 => X"000000fa",
    1752 => X"00000000",
    1753 => X"0000d1b7",
    1754 => X"00000ddb",
    1755 => X"000000fa",
    1756 => X"00000000",
    1757 => X"0000d1b7",
    1758 => X"00000de0",
    1759 => X"000000fa",
    1760 => X"00000000",
    1761 => X"0000d1b7",
    1762 => X"00000de4",
    1763 => X"000000fa",
    1764 => X"00000000",
    1765 => X"0000d1b7",
    1766 => X"00000de8",
    1767 => X"000000fa",
    1768 => X"00000000",
    1769 => X"0000d1b7",
    1770 => X"00000dec",
    1771 => X"000000fa",
    1772 => X"00000000",
    1773 => X"0000d1b7",
    1774 => X"00000df1",
    1775 => X"000000fa",
    1776 => X"00000000",
    1777 => X"0000d1b7",
    1778 => X"00000df5",
    1779 => X"000000fa",
    1780 => X"00000000",
    1781 => X"0000d1b7",
    1782 => X"00000df9",
    1783 => X"000000fa",
    1784 => X"00000000",
    1785 => X"0000d1b7",
    1786 => X"00000dfc",
    1787 => X"000000fa",
    1788 => X"00000000",
    1789 => X"0000d1b7",
    1790 => X"00000e00",
    1791 => X"000000fa",
    1792 => X"00000000",
    1793 => X"0000d1b7",
    1794 => X"00000e04",
    1795 => X"000000fa",
    1796 => X"00000000",
    1797 => X"0000d1b7",
    1798 => X"00000e08",
    1799 => X"000000fa",
    1800 => X"00000000",
    1801 => X"0000d1b7",
    1802 => X"00000e0b",
    1803 => X"000000fa",
    1804 => X"00000000",
    1805 => X"0000d1b7",
    1806 => X"00000e0f",
    1807 => X"000000fa",
    1808 => X"00000000",
    1809 => X"0000d1b7",
    1810 => X"00000e12",
    1811 => X"000000fa",
    1812 => X"00000000",
    1813 => X"0000d1b7",
    1814 => X"00000e16",
    1815 => X"000000fa",
    1816 => X"00000000",
    1817 => X"0000d1b7",
    1818 => X"00000e19",
    1819 => X"000000fa",
    1820 => X"00000000",
    1821 => X"0000d1b7",
    1822 => X"00000e1c",
    1823 => X"000000fa",
    1824 => X"00000000",
    1825 => X"0000d1b7",
    1826 => X"00000e20",
    1827 => X"000000fa",
    1828 => X"00000000",
    1829 => X"0000d1b7",
    1830 => X"00000e23",
    1831 => X"000000fa",
    1832 => X"00000000",
    1833 => X"0000d1b7",
    1834 => X"00000e26",
    1835 => X"000000fa",
    1836 => X"00000000",
    1837 => X"0000d1b7",
    1838 => X"00000e29",
    1839 => X"000000fa",
    1840 => X"00000000",
    1841 => X"0000d1b7",
    1842 => X"00000e2c",
    1843 => X"000000fa",
    1844 => X"00000000",
    1845 => X"0000d1b7",
    1846 => X"00000e2e",
    1847 => X"000000fa",
    1848 => X"00000000",
    1849 => X"0000d1b7",
    1850 => X"00000e31",
    1851 => X"000000fa",
    1852 => X"00000000",
    1853 => X"0000d1b7",
    1854 => X"00000e34",
    1855 => X"000000fa",
    1856 => X"00000000",
    1857 => X"0000d1b7",
    1858 => X"00000e37",
    1859 => X"000000fa",
    1860 => X"00000000",
    1861 => X"0000d1b7",
    1862 => X"00000e39",
    1863 => X"000000fa",
    1864 => X"00000000",
    1865 => X"0000d1b7",
    1866 => X"00000e3c",
    1867 => X"000000fa",
    1868 => X"00000000",
    1869 => X"0000d1b7",
    1870 => X"00000e3e",
    1871 => X"000000fa",
    1872 => X"00000000",
    1873 => X"0000d1b7",
    1874 => X"00000e40",
    1875 => X"000000fa",
    1876 => X"00000000",
    1877 => X"0000d1b7",
    1878 => X"00000e43",
    1879 => X"000000fa",
    1880 => X"00000000",
    1881 => X"0000d1b7",
    1882 => X"00000e45",
    1883 => X"000000fa",
    1884 => X"00000000",
    1885 => X"0000d1b7",
    1886 => X"00000e47",
    1887 => X"000000fa",
    1888 => X"00000000",
    1889 => X"0000d1b7",
    1890 => X"00000e49",
    1891 => X"000000fa",
    1892 => X"00000000",
    1893 => X"0000d1b7",
    1894 => X"00000e4b",
    1895 => X"000000fa",
    1896 => X"00000000",
    1897 => X"0000d1b7",
    1898 => X"00000e4d",
    1899 => X"000000fa",
    1900 => X"00000000",
    1901 => X"0000d1b7",
    1902 => X"00000e4f",
    1903 => X"000000fa",
    1904 => X"00000000",
    1905 => X"0000d1b7",
    1906 => X"00000e51",
    1907 => X"000000fa",
    1908 => X"00000000",
    1909 => X"0000d1b7",
    1910 => X"00000e52",
    1911 => X"000000fa",
    1912 => X"00000000",
    1913 => X"0000d1b7",
    1914 => X"00000e54",
    1915 => X"000000fa",
    1916 => X"00000000",
    1917 => X"0000d1b7",
    1918 => X"00000e55",
    1919 => X"000000fa",
    1920 => X"00000000",
    1921 => X"0000d1b7",
    1922 => X"00000e57",
    1923 => X"000000fa",
    1924 => X"00000000",
    1925 => X"0000d1b7",
    1926 => X"00000e58",
    1927 => X"000000fa",
    1928 => X"00000000",
    1929 => X"0000d1b7",
    1930 => X"00000e5a",
    1931 => X"000000fa",
    1932 => X"00000000",
    1933 => X"0000d1b7",
    1934 => X"00000e5b",
    1935 => X"000000fa",
    1936 => X"00000000",
    1937 => X"0000d1b7",
    1938 => X"00000e5c",
    1939 => X"000000fa",
    1940 => X"00000000",
    1941 => X"0000d1b7",
    1942 => X"00000e5d",
    1943 => X"000000fa",
    1944 => X"00000000",
    1945 => X"0000d1b7",
    1946 => X"00000e5e",
    1947 => X"000000fa",
    1948 => X"00000000",
    1949 => X"0000d1b7",
    1950 => X"00000e5f",
    1951 => X"000000fa",
    1952 => X"00000000",
    1953 => X"0000d1b7",
    1954 => X"00000e60",
    1955 => X"000000fa",
    1956 => X"00000000",
    1957 => X"0000d1b7",
    1958 => X"00000e61",
    1959 => X"000000fa",
    1960 => X"00000000",
    1961 => X"0000d1b7",
    1962 => X"00000e62",
    1963 => X"000000fa",
    1964 => X"00000000",
    1965 => X"0000d1b7",
    1966 => X"00000e63",
    1967 => X"000000fa",
    1968 => X"00000000",
    1969 => X"0000d1b7",
    1970 => X"00000e63",
    1971 => X"000000fa",
    1972 => X"00000000",
    1973 => X"0000d1b7",
    1974 => X"00000e64",
    1975 => X"000000fa",
    1976 => X"00000000",
    1977 => X"0000d1b7",
    1978 => X"00000e64",
    1979 => X"000000fa",
    1980 => X"00000000",
    1981 => X"0000d1b7",
    1982 => X"00000e65",
    1983 => X"000000fa",
    1984 => X"00000000",
    1985 => X"0000d1b7",
    1986 => X"00000e65",
    1987 => X"000000fa",
    1988 => X"00000000",
    1989 => X"0000d1b7",
    1990 => X"00000e65",
    1991 => X"000000fa",
    1992 => X"00000000",
    1993 => X"0000d1b7",
    1994 => X"00000e65",
    1995 => X"000000fa",
    1996 => X"00000000",
    1997 => X"0000d1b7",
    1998 => X"00000e65",
    1999 => X"000000fa",
    2000 => X"00000000",
    2001 => X"0000d1b7",
    2002 => X"00000e66",
    2003 => X"000000fa",
    2004 => X"00000000",
    2005 => X"0000d1b7",
    2006 => X"00000e65",
    2007 => X"000000fa",
    2008 => X"00000000",
    2009 => X"0000d1b7",
    2010 => X"00000e65",
    2011 => X"000000fa",
    2012 => X"00000000",
    2013 => X"0000d1b7",
    2014 => X"00000e65",
    2015 => X"000000fa",
    2016 => X"00000000",
    2017 => X"0000d1b7",
    2018 => X"00000e65",
    2019 => X"000000fa",
    2020 => X"00000000",
    2021 => X"0000d1b7",
    2022 => X"00000e65",
    2023 => X"000000fa",
    2024 => X"00000000",
    2025 => X"0000d1b7",
    2026 => X"00000e64",
    2027 => X"000000fa",
    2028 => X"00000000",
    2029 => X"0000d1b7",
    2030 => X"00000e64",
    2031 => X"000000fa",
    2032 => X"00000000",
    2033 => X"0000d1b7",
    2034 => X"00000e63",
    2035 => X"000000fa",
    2036 => X"00000000",
    2037 => X"0000d1b7",
    2038 => X"00000e63",
    2039 => X"000000fa",
    2040 => X"00000000",
    2041 => X"0000d1b7",
    2042 => X"00000e62",
    2043 => X"000000fa",
    2044 => X"00000000",
    2045 => X"0000d1b7",
    2046 => X"00000e61",
    2047 => X"000000fa",
    2048 => X"00000000",
    2049 => X"0000d1b7",
    2050 => X"00000e60",
    2051 => X"000000fa",
    2052 => X"00000000",
    2053 => X"0000d1b7",
    2054 => X"00000e5f",
    2055 => X"000000fa",
    2056 => X"00000000",
    2057 => X"0000d1b7",
    2058 => X"00000e5e",
    2059 => X"000000fa",
    2060 => X"00000000",
    2061 => X"0000d1b7",
    2062 => X"00000e5d",
    2063 => X"000000fa",
    2064 => X"00000000",
    2065 => X"0000d1b7",
    2066 => X"00000e5c",
    2067 => X"000000fa",
    2068 => X"00000000",
    2069 => X"0000d1b7",
    2070 => X"00000e5b",
    2071 => X"000000fa",
    2072 => X"00000000",
    2073 => X"0000d1b7",
    2074 => X"00000e5a",
    2075 => X"000000fa",
    2076 => X"00000000",
    2077 => X"0000d1b7",
    2078 => X"00000e58",
    2079 => X"000000fa",
    2080 => X"00000000",
    2081 => X"0000d1b7",
    2082 => X"00000e57",
    2083 => X"000000fa",
    2084 => X"00000000",
    2085 => X"0000d1b7",
    2086 => X"00000e55",
    2087 => X"000000fa",
    2088 => X"00000000",
    2089 => X"0000d1b7",
    2090 => X"00000e54",
    2091 => X"000000fa",
    2092 => X"00000000",
    2093 => X"0000d1b7",
    2094 => X"00000e52",
    2095 => X"000000fa",
    2096 => X"00000000",
    2097 => X"0000d1b7",
    2098 => X"00000e51",
    2099 => X"000000fa",
    2100 => X"00000000",
    2101 => X"0000d1b7",
    2102 => X"00000e4f",
    2103 => X"000000fa",
    2104 => X"00000000",
    2105 => X"0000d1b7",
    2106 => X"00000e4d",
    2107 => X"000000fa",
    2108 => X"00000000",
    2109 => X"0000d1b7",
    2110 => X"00000e4b",
    2111 => X"000000fa",
    2112 => X"00000000",
    2113 => X"0000d1b7",
    2114 => X"00000e49",
    2115 => X"000000fa",
    2116 => X"00000000",
    2117 => X"0000d1b7",
    2118 => X"00000e47",
    2119 => X"000000fa",
    2120 => X"00000000",
    2121 => X"0000d1b7",
    2122 => X"00000e45",
    2123 => X"000000fa",
    2124 => X"00000000",
    2125 => X"0000d1b7",
    2126 => X"00000e43",
    2127 => X"000000fa",
    2128 => X"00000000",
    2129 => X"0000d1b7",
    2130 => X"00000e40",
    2131 => X"000000fa",
    2132 => X"00000000",
    2133 => X"0000d1b7",
    2134 => X"00000e3e",
    2135 => X"000000fa",
    2136 => X"00000000",
    2137 => X"0000d1b7",
    2138 => X"00000e3c",
    2139 => X"000000fa",
    2140 => X"00000000",
    2141 => X"0000d1b7",
    2142 => X"00000e39",
    2143 => X"000000fa",
    2144 => X"00000000",
    2145 => X"0000d1b7",
    2146 => X"00000e37",
    2147 => X"000000fa",
    2148 => X"00000000",
    2149 => X"0000d1b7",
    2150 => X"00000e34",
    2151 => X"000000fa",
    2152 => X"00000000",
    2153 => X"0000d1b7",
    2154 => X"00000e31",
    2155 => X"000000fa",
    2156 => X"00000000",
    2157 => X"0000d1b7",
    2158 => X"00000e2e",
    2159 => X"000000fa",
    2160 => X"00000000",
    2161 => X"0000d1b7",
    2162 => X"00000e2c",
    2163 => X"000000fa",
    2164 => X"00000000",
    2165 => X"0000d1b7",
    2166 => X"00000e29",
    2167 => X"000000fa",
    2168 => X"00000000",
    2169 => X"0000d1b7",
    2170 => X"00000e26",
    2171 => X"000000fa",
    2172 => X"00000000",
    2173 => X"0000d1b7",
    2174 => X"00000e23",
    2175 => X"000000fa",
    2176 => X"00000000",
    2177 => X"0000d1b7",
    2178 => X"00000e20",
    2179 => X"000000fa",
    2180 => X"00000000",
    2181 => X"0000d1b7",
    2182 => X"00000e1c",
    2183 => X"000000fa",
    2184 => X"00000000",
    2185 => X"0000d1b7",
    2186 => X"00000e19",
    2187 => X"000000fa",
    2188 => X"00000000",
    2189 => X"0000d1b7",
    2190 => X"00000e16",
    2191 => X"000000fa",
    2192 => X"00000000",
    2193 => X"0000d1b7",
    2194 => X"00000e12",
    2195 => X"000000fa",
    2196 => X"00000000",
    2197 => X"0000d1b7",
    2198 => X"00000e0f",
    2199 => X"000000fa",
    2200 => X"00000000",
    2201 => X"0000d1b7",
    2202 => X"00000e0b",
    2203 => X"000000fa",
    2204 => X"00000000",
    2205 => X"0000d1b7",
    2206 => X"00000e08",
    2207 => X"000000fa",
    2208 => X"00000000",
    2209 => X"0000d1b7",
    2210 => X"00000e04",
    2211 => X"000000fa",
    2212 => X"00000000",
    2213 => X"0000d1b7",
    2214 => X"00000e00",
    2215 => X"000000fa",
    2216 => X"00000000",
    2217 => X"0000d1b7",
    2218 => X"00000dfc",
    2219 => X"000000fa",
    2220 => X"00000000",
    2221 => X"0000d1b7",
    2222 => X"00000df9",
    2223 => X"000000fa",
    2224 => X"00000000",
    2225 => X"0000d1b7",
    2226 => X"00000df5",
    2227 => X"000000fa",
    2228 => X"00000000",
    2229 => X"0000d1b7",
    2230 => X"00000df1",
    2231 => X"000000fa",
    2232 => X"00000000",
    2233 => X"0000d1b7",
    2234 => X"00000dec",
    2235 => X"000000fa",
    2236 => X"00000000",
    2237 => X"0000d1b7",
    2238 => X"00000de8",
    2239 => X"000000fa",
    2240 => X"00000000",
    2241 => X"0000d1b7",
    2242 => X"00000de4",
    2243 => X"000000fa",
    2244 => X"00000000",
    2245 => X"0000d1b7",
    2246 => X"00000de0",
    2247 => X"000000fa",
    2248 => X"00000000",
    2249 => X"0000d1b7",
    2250 => X"00000ddb",
    2251 => X"000000fa",
    2252 => X"00000000",
    2253 => X"0000d1b7",
    2254 => X"00000dd7",
    2255 => X"000000fa",
    2256 => X"00000000",
    2257 => X"0000d1b7",
    2258 => X"00000dd3",
    2259 => X"000000fa",
    2260 => X"00000000",
    2261 => X"0000d1b7",
    2262 => X"00000dce",
    2263 => X"000000fa",
    2264 => X"00000000",
    2265 => X"0000d1b7",
    2266 => X"00000dc9",
    2267 => X"000000fa",
    2268 => X"00000000",
    2269 => X"0000d1b7",
    2270 => X"00000dc5",
    2271 => X"000000fa",
    2272 => X"00000000",
    2273 => X"0000d1b7",
    2274 => X"00000dc0",
    2275 => X"000000fa",
    2276 => X"00000000",
    2277 => X"0000d1b7",
    2278 => X"00000dbb",
    2279 => X"000000fa",
    2280 => X"00000000",
    2281 => X"0000d1b7",
    2282 => X"00000db6",
    2283 => X"000000fa",
    2284 => X"00000000",
    2285 => X"0000d1b7",
    2286 => X"00000db1",
    2287 => X"000000fa",
    2288 => X"00000000",
    2289 => X"0000d1b7",
    2290 => X"00000dac",
    2291 => X"000000fa",
    2292 => X"00000000",
    2293 => X"0000d1b7",
    2294 => X"00000da7",
    2295 => X"000000fa",
    2296 => X"00000000",
    2297 => X"0000d1b7",
    2298 => X"00000da2",
    2299 => X"000000fa",
    2300 => X"00000000",
    2301 => X"0000d1b7",
    2302 => X"00000d9d",
    2303 => X"000000fa",
    2304 => X"00000000",
    2305 => X"0000d1b7",
    2306 => X"00000d97",
    2307 => X"000000fa",
    2308 => X"00000000",
    2309 => X"0000d1b7",
    2310 => X"00000d92",
    2311 => X"000000fa",
    2312 => X"00000000",
    2313 => X"0000d1b7",
    2314 => X"00000d8d",
    2315 => X"000000fa",
    2316 => X"00000000",
    2317 => X"0000d1b7",
    2318 => X"00000d87",
    2319 => X"000000fa",
    2320 => X"00000000",
    2321 => X"0000d1b7",
    2322 => X"00000d82",
    2323 => X"000000fa",
    2324 => X"00000000",
    2325 => X"0000d1b7",
    2326 => X"00000d7c",
    2327 => X"000000fa",
    2328 => X"00000000",
    2329 => X"0000d1b7",
    2330 => X"00000d76",
    2331 => X"000000fa",
    2332 => X"00000000",
    2333 => X"0000d1b7",
    2334 => X"00000d71",
    2335 => X"000000fa",
    2336 => X"00000000",
    2337 => X"0000d1b7",
    2338 => X"00000d6b",
    2339 => X"000000fa",
    2340 => X"00000000",
    2341 => X"0000d1b7",
    2342 => X"00000d65",
    2343 => X"000000fa",
    2344 => X"00000000",
    2345 => X"0000d1b7",
    2346 => X"00000d5f",
    2347 => X"000000fa",
    2348 => X"00000000",
    2349 => X"0000d1b7",
    2350 => X"00000d59",
    2351 => X"000000fa",
    2352 => X"00000000",
    2353 => X"0000d1b7",
    2354 => X"00000d53",
    2355 => X"000000fa",
    2356 => X"00000000",
    2357 => X"0000d1b7",
    2358 => X"00000d4d",
    2359 => X"000000fa",
    2360 => X"00000000",
    2361 => X"0000d1b7",
    2362 => X"00000d47",
    2363 => X"000000fa",
    2364 => X"00000000",
    2365 => X"0000d1b7",
    2366 => X"00000d40",
    2367 => X"000000fa",
    2368 => X"00000000",
    2369 => X"0000d1b7",
    2370 => X"00000d3a",
    2371 => X"000000fa",
    2372 => X"00000000",
    2373 => X"0000d1b7",
    2374 => X"00000d34",
    2375 => X"000000fa",
    2376 => X"00000000",
    2377 => X"0000d1b7",
    2378 => X"00000d2d",
    2379 => X"000000fa",
    2380 => X"00000000",
    2381 => X"0000d1b7",
    2382 => X"00000d27",
    2383 => X"000000fa",
    2384 => X"00000000",
    2385 => X"0000d1b7",
    2386 => X"00000d20",
    2387 => X"000000fa",
    2388 => X"00000000",
    2389 => X"0000d1b7",
    2390 => X"00000d1a",
    2391 => X"000000fa",
    2392 => X"00000000",
    2393 => X"0000d1b7",
    2394 => X"00000d13",
    2395 => X"000000fa",
    2396 => X"00000000",
    2397 => X"0000d1b7",
    2398 => X"00000d0c",
    2399 => X"000000fa",
    2400 => X"00000000",
    2401 => X"0000d1b7",
    2402 => X"00000d06",
    2403 => X"000000fa",
    2404 => X"00000000",
    2405 => X"0000d1b7",
    2406 => X"00000cff",
    2407 => X"000000fa",
    2408 => X"00000000",
    2409 => X"0000d1b7",
    2410 => X"00000cf8",
    2411 => X"000000fa",
    2412 => X"00000000",
    2413 => X"0000d1b7",
    2414 => X"00000cf1",
    2415 => X"000000fa",
    2416 => X"00000000",
    2417 => X"0000d1b7",
    2418 => X"00000cea",
    2419 => X"000000fa",
    2420 => X"00000000",
    2421 => X"0000d1b7",
    2422 => X"00000ce3",
    2423 => X"000000fa",
    2424 => X"00000000",
    2425 => X"0000d1b7",
    2426 => X"00000cdc",
    2427 => X"000000fa",
    2428 => X"00000000",
    2429 => X"0000d1b7",
    2430 => X"00000cd5",
    2431 => X"000000fa",
    2432 => X"00000000",
    2433 => X"0000d1b7",
    2434 => X"00000ccd",
    2435 => X"000000fa",
    2436 => X"00000000",
    2437 => X"0000d1b7",
    2438 => X"00000cc6",
    2439 => X"000000fa",
    2440 => X"00000000",
    2441 => X"0000d1b7",
    2442 => X"00000cbf",
    2443 => X"000000fa",
    2444 => X"00000000",
    2445 => X"0000d1b7",
    2446 => X"00000cb7",
    2447 => X"000000fa",
    2448 => X"00000000",
    2449 => X"0000d1b7",
    2450 => X"00000cb0",
    2451 => X"000000fa",
    2452 => X"00000000",
    2453 => X"0000d1b7",
    2454 => X"00000ca8",
    2455 => X"000000fa",
    2456 => X"00000000",
    2457 => X"0000d1b7",
    2458 => X"00000ca1",
    2459 => X"000000fa",
    2460 => X"00000000",
    2461 => X"0000d1b7",
    2462 => X"00000c99",
    2463 => X"000000fa",
    2464 => X"00000000",
    2465 => X"0000d1b7",
    2466 => X"00000c91",
    2467 => X"000000fa",
    2468 => X"00000000",
    2469 => X"0000d1b7",
    2470 => X"00000c8a",
    2471 => X"000000fa",
    2472 => X"00000000",
    2473 => X"0000d1b7",
    2474 => X"00000c82",
    2475 => X"000000fa",
    2476 => X"00000000",
    2477 => X"0000d1b7",
    2478 => X"00000c7a",
    2479 => X"000000fa",
    2480 => X"00000000",
    2481 => X"0000d1b7",
    2482 => X"00000c72",
    2483 => X"000000fa",
    2484 => X"00000000",
    2485 => X"0000d1b7",
    2486 => X"00000c6a",
    2487 => X"000000fa",
    2488 => X"00000000",
    2489 => X"0000d1b7",
    2490 => X"00000c62",
    2491 => X"000000fa",
    2492 => X"00000000",
    2493 => X"0000d1b7",
    2494 => X"00000c5a",
    2495 => X"000000fa",
    2496 => X"00000000",
    2497 => X"0000d1b7",
    2498 => X"00000c52",
    2499 => X"000000fa",
    2500 => X"00000000",
    2501 => X"0000d1b7",
    2502 => X"00000c4a",
    2503 => X"000000fa",
    2504 => X"00000000",
    2505 => X"0000d1b7",
    2506 => X"00000c42",
    2507 => X"000000fa",
    2508 => X"00000000",
    2509 => X"0000d1b7",
    2510 => X"00000c39",
    2511 => X"000000fa",
    2512 => X"00000000",
    2513 => X"0000d1b7",
    2514 => X"00000c31",
    2515 => X"000000fa",
    2516 => X"00000000",
    2517 => X"0000d1b7",
    2518 => X"00000c29",
    2519 => X"000000fa",
    2520 => X"00000000",
    2521 => X"0000d1b7",
    2522 => X"00000c20",
    2523 => X"000000fa",
    2524 => X"00000000",
    2525 => X"0000d1b7",
    2526 => X"00000c18",
    2527 => X"000000fa",
    2528 => X"00000000",
    2529 => X"0000d1b7",
    2530 => X"00000c0f",
    2531 => X"000000fa",
    2532 => X"00000000",
    2533 => X"0000d1b7",
    2534 => X"00000c07",
    2535 => X"000000fa",
    2536 => X"00000000",
    2537 => X"0000d1b7",
    2538 => X"00000bfe",
    2539 => X"000000fa",
    2540 => X"00000000",
    2541 => X"0000d1b7",
    2542 => X"00000bf5",
    2543 => X"000000fa",
    2544 => X"00000000",
    2545 => X"0000d1b7",
    2546 => X"00000bed",
    2547 => X"000000fa",
    2548 => X"00000000",
    2549 => X"0000d1b7",
    2550 => X"00000be4",
    2551 => X"000000fa",
    2552 => X"00000000",
    2553 => X"0000d1b7",
    2554 => X"00000bdb",
    2555 => X"000000fa",
    2556 => X"00000000",
    2557 => X"0000d1b7",
    2558 => X"00000bd2",
    2559 => X"000000fa",
    2560 => X"00000000",
    2561 => X"0000d1b7",
    2562 => X"00000bc9",
    2563 => X"000000fa",
    2564 => X"00000000",
    2565 => X"0000d1b7",
    2566 => X"00000bc0",
    2567 => X"000000fa",
    2568 => X"00000000",
    2569 => X"0000d1b7",
    2570 => X"00000bb7",
    2571 => X"000000fa",
    2572 => X"00000000",
    2573 => X"0000d1b7",
    2574 => X"00000bae",
    2575 => X"000000fa",
    2576 => X"00000000",
    2577 => X"0000d1b7",
    2578 => X"00000ba5",
    2579 => X"000000fa",
    2580 => X"00000000",
    2581 => X"0000d1b7",
    2582 => X"00000b9c",
    2583 => X"000000fa",
    2584 => X"00000000",
    2585 => X"0000d1b7",
    2586 => X"00000b93",
    2587 => X"000000fa",
    2588 => X"00000000",
    2589 => X"0000d1b7",
    2590 => X"00000b8a",
    2591 => X"000000fa",
    2592 => X"00000000",
    2593 => X"0000d1b7",
    2594 => X"00000b81",
    2595 => X"000000fa",
    2596 => X"00000000",
    2597 => X"0000d1b7",
    2598 => X"00000b77",
    2599 => X"000000fa",
    2600 => X"00000000",
    2601 => X"0000d1b7",
    2602 => X"00000b6e",
    2603 => X"000000fa",
    2604 => X"00000000",
    2605 => X"0000d1b7",
    2606 => X"00000b65",
    2607 => X"000000fa",
    2608 => X"00000000",
    2609 => X"0000d1b7",
    2610 => X"00000b5b",
    2611 => X"000000fa",
    2612 => X"00000000",
    2613 => X"0000d1b7",
    2614 => X"00000b52",
    2615 => X"000000fa",
    2616 => X"00000000",
    2617 => X"0000d1b7",
    2618 => X"00000b48",
    2619 => X"000000fa",
    2620 => X"00000000",
    2621 => X"0000d1b7",
    2622 => X"00000b3f",
    2623 => X"000000fa",
    2624 => X"00000000",
    2625 => X"0000d1b7",
    2626 => X"00000b35",
    2627 => X"000000fa",
    2628 => X"00000000",
    2629 => X"0000d1b7",
    2630 => X"00000b2b",
    2631 => X"000000fa",
    2632 => X"00000000",
    2633 => X"0000d1b7",
    2634 => X"00000b22",
    2635 => X"000000fa",
    2636 => X"00000000",
    2637 => X"0000d1b7",
    2638 => X"00000b18",
    2639 => X"000000fa",
    2640 => X"00000000",
    2641 => X"0000d1b7",
    2642 => X"00000b0e",
    2643 => X"000000fa",
    2644 => X"00000000",
    2645 => X"0000d1b7",
    2646 => X"00000b04",
    2647 => X"000000fa",
    2648 => X"00000000",
    2649 => X"0000d1b7",
    2650 => X"00000afb",
    2651 => X"000000fa",
    2652 => X"00000000",
    2653 => X"0000d1b7",
    2654 => X"00000af1",
    2655 => X"000000fa",
    2656 => X"00000000",
    2657 => X"0000d1b7",
    2658 => X"00000ae7",
    2659 => X"000000fa",
    2660 => X"00000000",
    2661 => X"0000d1b7",
    2662 => X"00000add",
    2663 => X"000000fa",
    2664 => X"00000000",
    2665 => X"0000d1b7",
    2666 => X"00000ad3",
    2667 => X"000000fa",
    2668 => X"00000000",
    2669 => X"0000d1b7",
    2670 => X"00000ac9",
    2671 => X"000000fa",
    2672 => X"00000000",
    2673 => X"0000d1b7",
    2674 => X"00000abf",
    2675 => X"000000fa",
    2676 => X"00000000",
    2677 => X"0000d1b7",
    2678 => X"00000ab5",
    2679 => X"000000fa",
    2680 => X"00000000",
    2681 => X"0000d1b7",
    2682 => X"00000aab",
    2683 => X"000000fa",
    2684 => X"00000000",
    2685 => X"0000d1b7",
    2686 => X"00000aa0",
    2687 => X"000000fa",
    2688 => X"00000000",
    2689 => X"0000d1b7",
    2690 => X"00000a96",
    2691 => X"000000fa",
    2692 => X"00000000",
    2693 => X"0000d1b7",
    2694 => X"00000a8c",
    2695 => X"000000fa",
    2696 => X"00000000",
    2697 => X"0000d1b7",
    2698 => X"00000a82",
    2699 => X"000000fa",
    2700 => X"00000000",
    2701 => X"0000d1b7",
    2702 => X"00000a77",
    2703 => X"000000fa",
    2704 => X"00000000",
    2705 => X"0000d1b7",
    2706 => X"00000a6d",
    2707 => X"000000fa",
    2708 => X"00000000",
    2709 => X"0000d1b7",
    2710 => X"00000a63",
    2711 => X"000000fa",
    2712 => X"00000000",
    2713 => X"0000d1b7",
    2714 => X"00000a58",
    2715 => X"000000fa",
    2716 => X"00000000",
    2717 => X"0000d1b7",
    2718 => X"00000a4e",
    2719 => X"000000fa",
    2720 => X"00000000",
    2721 => X"0000d1b7",
    2722 => X"00000a43",
    2723 => X"000000fa",
    2724 => X"00000000",
    2725 => X"0000d1b7",
    2726 => X"00000a39",
    2727 => X"000000fa",
    2728 => X"00000000",
    2729 => X"0000d1b7",
    2730 => X"00000a2e",
    2731 => X"000000fa",
    2732 => X"00000000",
    2733 => X"0000d1b7",
    2734 => X"00000a24",
    2735 => X"000000fa",
    2736 => X"00000000",
    2737 => X"0000d1b7",
    2738 => X"00000a19",
    2739 => X"000000fa",
    2740 => X"00000000",
    2741 => X"0000d1b7",
    2742 => X"00000a0f",
    2743 => X"000000fa",
    2744 => X"00000000",
    2745 => X"0000d1b7",
    2746 => X"00000a04",
    2747 => X"000000fa",
    2748 => X"00000000",
    2749 => X"0000d1b7",
    2750 => X"000009f9",
    2751 => X"000000fa",
    2752 => X"00000000",
    2753 => X"0000d1b7",
    2754 => X"000009ef",
    2755 => X"000000fa",
    2756 => X"00000000",
    2757 => X"0000d1b7",
    2758 => X"000009e4",
    2759 => X"000000fa",
    2760 => X"00000000",
    2761 => X"0000d1b7",
    2762 => X"000009d9",
    2763 => X"000000fa",
    2764 => X"00000000",
    2765 => X"0000d1b7",
    2766 => X"000009ce",
    2767 => X"000000fa",
    2768 => X"00000000",
    2769 => X"0000d1b7",
    2770 => X"000009c4",
    2771 => X"000000fa",
    2772 => X"00000000",
    2773 => X"0000d1b7",
    2774 => X"000009b9",
    2775 => X"000000fa",
    2776 => X"00000000",
    2777 => X"0000d1b7",
    2778 => X"000009ae",
    2779 => X"000000fa",
    2780 => X"00000000",
    2781 => X"0000d1b7",
    2782 => X"000009a3",
    2783 => X"000000fa",
    2784 => X"00000000",
    2785 => X"0000d1b7",
    2786 => X"00000998",
    2787 => X"000000fa",
    2788 => X"00000000",
    2789 => X"0000d1b7",
    2790 => X"0000098d",
    2791 => X"000000fa",
    2792 => X"00000000",
    2793 => X"0000d1b7",
    2794 => X"00000982",
    2795 => X"000000fa",
    2796 => X"00000000",
    2797 => X"0000d1b7",
    2798 => X"00000977",
    2799 => X"000000fa",
    2800 => X"00000000",
    2801 => X"0000d1b7",
    2802 => X"0000096c",
    2803 => X"000000fa",
    2804 => X"00000000",
    2805 => X"0000d1b7",
    2806 => X"00000961",
    2807 => X"000000fa",
    2808 => X"00000000",
    2809 => X"0000d1b7",
    2810 => X"00000956",
    2811 => X"000000fa",
    2812 => X"00000000",
    2813 => X"0000d1b7",
    2814 => X"0000094b",
    2815 => X"000000fa",
    2816 => X"00000000",
    2817 => X"0000d1b7",
    2818 => X"00000940",
    2819 => X"000000fa",
    2820 => X"00000000",
    2821 => X"0000d1b7",
    2822 => X"00000935",
    2823 => X"000000fa",
    2824 => X"00000000",
    2825 => X"0000d1b7",
    2826 => X"0000092a",
    2827 => X"000000fa",
    2828 => X"00000000",
    2829 => X"0000d1b7",
    2830 => X"0000091f",
    2831 => X"000000fa",
    2832 => X"00000000",
    2833 => X"0000d1b7",
    2834 => X"00000913",
    2835 => X"000000fa",
    2836 => X"00000000",
    2837 => X"0000d1b7",
    2838 => X"00000908",
    2839 => X"000000fa",
    2840 => X"00000000",
    2841 => X"0000d1b7",
    2842 => X"000008fd",
    2843 => X"000000fa",
    2844 => X"00000000",
    2845 => X"0000d1b7",
    2846 => X"000008f2",
    2847 => X"000000fa",
    2848 => X"00000000",
    2849 => X"0000d1b7",
    2850 => X"000008e7",
    2851 => X"000000fa",
    2852 => X"00000000",
    2853 => X"0000d1b7",
    2854 => X"000008db",
    2855 => X"000000fa",
    2856 => X"00000000",
    2857 => X"0000d1b7",
    2858 => X"000008d0",
    2859 => X"000000fa",
    2860 => X"00000000",
    2861 => X"0000d1b7",
    2862 => X"000008c5",
    2863 => X"000000fa",
    2864 => X"00000000",
    2865 => X"0000d1b7",
    2866 => X"000008b9",
    2867 => X"000000fa",
    2868 => X"00000000",
    2869 => X"0000d1b7",
    2870 => X"000008ae",
    2871 => X"000000fa",
    2872 => X"00000000",
    2873 => X"0000d1b7",
    2874 => X"000008a3",
    2875 => X"000000fa",
    2876 => X"00000000",
    2877 => X"0000d1b7",
    2878 => X"00000897",
    2879 => X"000000fa",
    2880 => X"00000000",
    2881 => X"0000d1b7",
    2882 => X"0000088c",
    2883 => X"000000fa",
    2884 => X"00000000",
    2885 => X"0000d1b7",
    2886 => X"00000881",
    2887 => X"000000fa",
    2888 => X"00000000",
    2889 => X"0000d1b7",
    2890 => X"00000875",
    2891 => X"000000fa",
    2892 => X"00000000",
    2893 => X"0000d1b7",
    2894 => X"0000086a",
    2895 => X"000000fa",
    2896 => X"00000000",
    2897 => X"0000d1b7",
    2898 => X"0000085e",
    2899 => X"000000fa",
    2900 => X"00000000",
    2901 => X"0000d1b7",
    2902 => X"00000853",
    2903 => X"000000fa",
    2904 => X"00000000",
    2905 => X"0000d1b7",
    2906 => X"00000848",
    2907 => X"000000fa",
    2908 => X"00000000",
    2909 => X"0000d1b7",
    2910 => X"0000083c",
    2911 => X"000000fa",
    2912 => X"00000000",
    2913 => X"0000d1b7",
    2914 => X"00000831",
    2915 => X"000000fa",
    2916 => X"00000000",
    2917 => X"0000d1b7",
    2918 => X"00000825",
    2919 => X"000000fa",
    2920 => X"00000000",
    2921 => X"0000d1b7",
    2922 => X"0000081a",
    2923 => X"000000fa",
    2924 => X"00000000",
    2925 => X"0000d1b7",
    2926 => X"0000080e",
    2927 => X"000000fa",
    2928 => X"00000000",
    2929 => X"0000d1b7",
    2930 => X"00000803",
    2931 => X"000000fa",
    2932 => X"00000000",
    2933 => X"0000d1b7",
    2934 => X"000007f7",
    2935 => X"000000fa",
    2936 => X"00000000",
    2937 => X"0000d1b7",
    2938 => X"000007ec",
    2939 => X"000000fa",
    2940 => X"00000000",
    2941 => X"0000d1b7",
    2942 => X"000007e0",
    2943 => X"000000fa",
    2944 => X"00000000",
    2945 => X"0000d1b7",
    2946 => X"000007d5",
    2947 => X"000000fa",
    2948 => X"00000000",
    2949 => X"0000d1b7",
    2950 => X"000007c9",
    2951 => X"000000fa",
    2952 => X"00000000",
    2953 => X"0000d1b7",
    2954 => X"000007be",
    2955 => X"000000fa",
    2956 => X"00000000",
    2957 => X"0000d1b7",
    2958 => X"000007b2",
    2959 => X"000000fa",
    2960 => X"00000000",
    2961 => X"0000d1b7",
    2962 => X"000007a6",
    2963 => X"000000fa",
    2964 => X"00000000",
    2965 => X"0000d1b7",
    2966 => X"0000079b",
    2967 => X"000000fa",
    2968 => X"00000000",
    2969 => X"0000d1b7",
    2970 => X"0000078f",
    2971 => X"000000fa",
    2972 => X"00000000",
    2973 => X"0000d1b7",
    2974 => X"00000784",
    2975 => X"000000fa",
    2976 => X"00000000",
    2977 => X"0000d1b7",
    2978 => X"00000778",
    2979 => X"000000fa",
    2980 => X"00000000",
    2981 => X"0000d1b7",
    2982 => X"0000076d",
    2983 => X"000000fa",
    2984 => X"00000000",
    2985 => X"0000d1b7",
    2986 => X"00000761",
    2987 => X"000000fa",
    2988 => X"00000000",
    2989 => X"0000d1b7",
    2990 => X"00000755",
    2991 => X"000000fa",
    2992 => X"00000000",
    2993 => X"0000d1b7",
    2994 => X"0000074a",
    2995 => X"000000fa",
    2996 => X"00000000",
    2997 => X"0000d1b7",
    2998 => X"0000073e",
    2999 => X"000000fa",
    3000 => X"00000000",
    3001 => X"0000d1b7",
    3002 => X"00000733",
    3003 => X"000000fa",
    3004 => X"00000000",
    3005 => X"0000d1b7",
    3006 => X"00000727",
    3007 => X"000000fa",
    3008 => X"00000000",
    3009 => X"0000d1b7",
    3010 => X"0000071c",
    3011 => X"000000fa",
    3012 => X"00000000",
    3013 => X"0000d1b7",
    3014 => X"00000710",
    3015 => X"000000fa",
    3016 => X"00000000",
    3017 => X"0000d1b7",
    3018 => X"00000704",
    3019 => X"000000fa",
    3020 => X"00000000",
    3021 => X"0000d1b7",
    3022 => X"000006f9",
    3023 => X"000000fa",
    3024 => X"00000000",
    3025 => X"0000d1b7",
    3026 => X"000006ed",
    3027 => X"000000fa",
    3028 => X"00000000",
    3029 => X"0000d1b7",
    3030 => X"000006e2",
    3031 => X"000000fa",
    3032 => X"00000000",
    3033 => X"0000d1b7",
    3034 => X"000006d6",
    3035 => X"000000fa",
    3036 => X"00000000",
    3037 => X"0000d1b7",
    3038 => X"000006cb",
    3039 => X"000000fa",
    3040 => X"00000000",
    3041 => X"0000d1b7",
    3042 => X"000006bf",
    3043 => X"000000fa",
    3044 => X"00000000",
    3045 => X"0000d1b7",
    3046 => X"000006b3",
    3047 => X"000000fa",
    3048 => X"00000000",
    3049 => X"0000d1b7",
    3050 => X"000006a8",
    3051 => X"000000fa",
    3052 => X"00000000",
    3053 => X"0000d1b7",
    3054 => X"0000069c",
    3055 => X"000000fa",
    3056 => X"00000000",
    3057 => X"0000d1b7",
    3058 => X"00000691",
    3059 => X"000000fa",
    3060 => X"00000000",
    3061 => X"0000d1b7",
    3062 => X"00000685",
    3063 => X"000000fa",
    3064 => X"00000000",
    3065 => X"0000d1b7",
    3066 => X"0000067a",
    3067 => X"000000fa",
    3068 => X"00000000",
    3069 => X"0000d1b7",
    3070 => X"0000066e",
    3071 => X"000000fa",
    3072 => X"00000000",
    3073 => X"0000d1b7",
    3074 => X"00000663",
    3075 => X"000000fa",
    3076 => X"00000000",
    3077 => X"0000d1b7",
    3078 => X"00000657",
    3079 => X"000000fa",
    3080 => X"00000000",
    3081 => X"0000d1b7",
    3082 => X"0000064c",
    3083 => X"000000fa",
    3084 => X"00000000",
    3085 => X"0000d1b7",
    3086 => X"00000640",
    3087 => X"000000fa",
    3088 => X"00000000",
    3089 => X"0000d1b7",
    3090 => X"00000635",
    3091 => X"000000fa",
    3092 => X"00000000",
    3093 => X"0000d1b7",
    3094 => X"00000629",
    3095 => X"000000fa",
    3096 => X"00000000",
    3097 => X"0000d1b7",
    3098 => X"0000061e",
    3099 => X"000000fa",
    3100 => X"00000000",
    3101 => X"0000d1b7",
    3102 => X"00000612",
    3103 => X"000000fa",
    3104 => X"00000000",
    3105 => X"0000d1b7",
    3106 => X"00000607",
    3107 => X"000000fa",
    3108 => X"00000000",
    3109 => X"0000d1b7",
    3110 => X"000005fc",
    3111 => X"000000fa",
    3112 => X"00000000",
    3113 => X"0000d1b7",
    3114 => X"000005f0",
    3115 => X"000000fa",
    3116 => X"00000000",
    3117 => X"0000d1b7",
    3118 => X"000005e5",
    3119 => X"000000fa",
    3120 => X"00000000",
    3121 => X"0000d1b7",
    3122 => X"000005d9",
    3123 => X"000000fa",
    3124 => X"00000000",
    3125 => X"0000d1b7",
    3126 => X"000005ce",
    3127 => X"000000fa",
    3128 => X"00000000",
    3129 => X"0000d1b7",
    3130 => X"000005c3",
    3131 => X"000000fa",
    3132 => X"00000000",
    3133 => X"0000d1b7",
    3134 => X"000005b7",
    3135 => X"000000fa",
    3136 => X"00000000",
    3137 => X"0000d1b7",
    3138 => X"000005ac",
    3139 => X"000000fa",
    3140 => X"00000000",
    3141 => X"0000d1b7",
    3142 => X"000005a1",
    3143 => X"000000fa",
    3144 => X"00000000",
    3145 => X"0000d1b7",
    3146 => X"00000595",
    3147 => X"000000fa",
    3148 => X"00000000",
    3149 => X"0000d1b7",
    3150 => X"0000058a",
    3151 => X"000000fa",
    3152 => X"00000000",
    3153 => X"0000d1b7",
    3154 => X"0000057f",
    3155 => X"000000fa",
    3156 => X"00000000",
    3157 => X"0000d1b7",
    3158 => X"00000574",
    3159 => X"000000fa",
    3160 => X"00000000",
    3161 => X"0000d1b7",
    3162 => X"00000568",
    3163 => X"000000fa",
    3164 => X"00000000",
    3165 => X"0000d1b7",
    3166 => X"0000055d",
    3167 => X"000000fa",
    3168 => X"00000000",
    3169 => X"0000d1b7",
    3170 => X"00000552",
    3171 => X"000000fa",
    3172 => X"00000000",
    3173 => X"0000d1b7",
    3174 => X"00000547",
    3175 => X"000000fa",
    3176 => X"00000000",
    3177 => X"0000d1b7",
    3178 => X"0000053c",
    3179 => X"000000fa",
    3180 => X"00000000",
    3181 => X"0000d1b7",
    3182 => X"00000531",
    3183 => X"000000fa",
    3184 => X"00000000",
    3185 => X"0000d1b7",
    3186 => X"00000526",
    3187 => X"000000fa",
    3188 => X"00000000",
    3189 => X"0000d1b7",
    3190 => X"0000051a",
    3191 => X"000000fa",
    3192 => X"00000000",
    3193 => X"0000d1b7",
    3194 => X"0000050f",
    3195 => X"000000fa",
    3196 => X"00000000",
    3197 => X"0000d1b7",
    3198 => X"00000504",
    3199 => X"000000fa",
    3200 => X"00000000",
    3201 => X"0000d1b7",
    3202 => X"000004f9",
    3203 => X"000000fa",
    3204 => X"00000000",
    3205 => X"0000d1b7",
    3206 => X"000004ee",
    3207 => X"000000fa",
    3208 => X"00000000",
    3209 => X"0000d1b7",
    3210 => X"000004e3",
    3211 => X"000000fa",
    3212 => X"00000000",
    3213 => X"0000d1b7",
    3214 => X"000004d8",
    3215 => X"000000fa",
    3216 => X"00000000",
    3217 => X"0000d1b7",
    3218 => X"000004cd",
    3219 => X"000000fa",
    3220 => X"00000000",
    3221 => X"0000d1b7",
    3222 => X"000004c3",
    3223 => X"000000fa",
    3224 => X"00000000",
    3225 => X"0000d1b7",
    3226 => X"000004b8",
    3227 => X"000000fa",
    3228 => X"00000000",
    3229 => X"0000d1b7",
    3230 => X"000004ad",
    3231 => X"000000fa",
    3232 => X"00000000",
    3233 => X"0000d1b7",
    3234 => X"000004a2",
    3235 => X"000000fa",
    3236 => X"00000000",
    3237 => X"0000d1b7",
    3238 => X"00000497",
    3239 => X"000000fa",
    3240 => X"00000000",
    3241 => X"0000d1b7",
    3242 => X"0000048c",
    3243 => X"000000fa",
    3244 => X"00000000",
    3245 => X"0000d1b7",
    3246 => X"00000482",
    3247 => X"000000fa",
    3248 => X"00000000",
    3249 => X"0000d1b7",
    3250 => X"00000477",
    3251 => X"000000fa",
    3252 => X"00000000",
    3253 => X"0000d1b7",
    3254 => X"0000046c",
    3255 => X"000000fa",
    3256 => X"00000000",
    3257 => X"0000d1b7",
    3258 => X"00000462",
    3259 => X"000000fa",
    3260 => X"00000000",
    3261 => X"0000d1b7",
    3262 => X"00000457",
    3263 => X"000000fa",
    3264 => X"00000000",
    3265 => X"0000d1b7",
    3266 => X"0000044c",
    3267 => X"000000fa",
    3268 => X"00000000",
    3269 => X"0000d1b7",
    3270 => X"00000442",
    3271 => X"000000fa",
    3272 => X"00000000",
    3273 => X"0000d1b7",
    3274 => X"00000437",
    3275 => X"000000fa",
    3276 => X"00000000",
    3277 => X"0000d1b7",
    3278 => X"0000042d",
    3279 => X"000000fa",
    3280 => X"00000000",
    3281 => X"0000d1b7",
    3282 => X"00000422",
    3283 => X"000000fa",
    3284 => X"00000000",
    3285 => X"0000d1b7",
    3286 => X"00000418",
    3287 => X"000000fa",
    3288 => X"00000000",
    3289 => X"0000d1b7",
    3290 => X"0000040d",
    3291 => X"000000fa",
    3292 => X"00000000",
    3293 => X"0000d1b7",
    3294 => X"00000403",
    3295 => X"000000fa",
    3296 => X"00000000",
    3297 => X"0000d1b7",
    3298 => X"000003f8",
    3299 => X"000000fa",
    3300 => X"00000000",
    3301 => X"0000d1b7",
    3302 => X"000003ee",
    3303 => X"000000fa",
    3304 => X"00000000",
    3305 => X"0000d1b7",
    3306 => X"000003e4",
    3307 => X"000000fa",
    3308 => X"00000000",
    3309 => X"0000d1b7",
    3310 => X"000003da",
    3311 => X"000000fa",
    3312 => X"00000000",
    3313 => X"0000d1b7",
    3314 => X"000003cf",
    3315 => X"000000fa",
    3316 => X"00000000",
    3317 => X"0000d1b7",
    3318 => X"000003c5",
    3319 => X"000000fa",
    3320 => X"00000000",
    3321 => X"0000d1b7",
    3322 => X"000003bb",
    3323 => X"000000fa",
    3324 => X"00000000",
    3325 => X"0000d1b7",
    3326 => X"000003b1",
    3327 => X"000000fa",
    3328 => X"00000000",
    3329 => X"0000d1b7",
    3330 => X"000003a7",
    3331 => X"000000fa",
    3332 => X"00000000",
    3333 => X"0000d1b7",
    3334 => X"0000039d",
    3335 => X"000000fa",
    3336 => X"00000000",
    3337 => X"0000d1b7",
    3338 => X"00000393",
    3339 => X"000000fa",
    3340 => X"00000000",
    3341 => X"0000d1b7",
    3342 => X"00000389",
    3343 => X"000000fa",
    3344 => X"00000000",
    3345 => X"0000d1b7",
    3346 => X"0000037f",
    3347 => X"000000fa",
    3348 => X"00000000",
    3349 => X"0000d1b7",
    3350 => X"00000375",
    3351 => X"000000fa",
    3352 => X"00000000",
    3353 => X"0000d1b7",
    3354 => X"0000036b",
    3355 => X"000000fa",
    3356 => X"00000000",
    3357 => X"0000d1b7",
    3358 => X"00000361",
    3359 => X"000000fa",
    3360 => X"00000000",
    3361 => X"0000d1b7",
    3362 => X"00000357",
    3363 => X"000000fa",
    3364 => X"00000000",
    3365 => X"0000d1b7",
    3366 => X"0000034e",
    3367 => X"000000fa",
    3368 => X"00000000",
    3369 => X"0000d1b7",
    3370 => X"00000344",
    3371 => X"000000fa",
    3372 => X"00000000",
    3373 => X"0000d1b7",
    3374 => X"0000033a",
    3375 => X"000000fa",
    3376 => X"00000000",
    3377 => X"0000d1b7",
    3378 => X"00000331",
    3379 => X"000000fa",
    3380 => X"00000000",
    3381 => X"0000d1b7",
    3382 => X"00000327",
    3383 => X"000000fa",
    3384 => X"00000000",
    3385 => X"0000d1b7",
    3386 => X"0000031d",
    3387 => X"000000fa",
    3388 => X"00000000",
    3389 => X"0000d1b7",
    3390 => X"00000314",
    3391 => X"000000fa",
    3392 => X"00000000",
    3393 => X"0000d1b7",
    3394 => X"0000030a",
    3395 => X"000000fa",
    3396 => X"00000000",
    3397 => X"0000d1b7",
    3398 => X"00000301",
    3399 => X"000000fa",
    3400 => X"00000000",
    3401 => X"0000d1b7",
    3402 => X"000002f8",
    3403 => X"000000fa",
    3404 => X"00000000",
    3405 => X"0000d1b7",
    3406 => X"000002ee",
    3407 => X"000000fa",
    3408 => X"00000000",
    3409 => X"0000d1b7",
    3410 => X"000002e5",
    3411 => X"000000fa",
    3412 => X"00000000",
    3413 => X"0000d1b7",
    3414 => X"000002dc",
    3415 => X"000000fa",
    3416 => X"00000000",
    3417 => X"0000d1b7",
    3418 => X"000002d2",
    3419 => X"000000fa",
    3420 => X"00000000",
    3421 => X"0000d1b7",
    3422 => X"000002c9",
    3423 => X"000000fa",
    3424 => X"00000000",
    3425 => X"0000d1b7",
    3426 => X"000002c0",
    3427 => X"000000fa",
    3428 => X"00000000",
    3429 => X"0000d1b7",
    3430 => X"000002b7",
    3431 => X"000000fa",
    3432 => X"00000000",
    3433 => X"0000d1b7",
    3434 => X"000002ae",
    3435 => X"000000fa",
    3436 => X"00000000",
    3437 => X"0000d1b7",
    3438 => X"000002a5",
    3439 => X"000000fa",
    3440 => X"00000000",
    3441 => X"0000d1b7",
    3442 => X"0000029c",
    3443 => X"000000fa",
    3444 => X"00000000",
    3445 => X"0000d1b7",
    3446 => X"00000293",
    3447 => X"000000fa",
    3448 => X"00000000",
    3449 => X"0000d1b7",
    3450 => X"0000028a",
    3451 => X"000000fa",
    3452 => X"00000000",
    3453 => X"0000d1b7",
    3454 => X"00000282",
    3455 => X"000000fa",
    3456 => X"00000000",
    3457 => X"0000d1b7",
    3458 => X"00000279",
    3459 => X"000000fa",
    3460 => X"00000000",
    3461 => X"0000d1b7",
    3462 => X"00000270",
    3463 => X"000000fa",
    3464 => X"00000000",
    3465 => X"0000d1b7",
    3466 => X"00000267",
    3467 => X"000000fa",
    3468 => X"00000000",
    3469 => X"0000d1b7",
    3470 => X"0000025f",
    3471 => X"000000fa",
    3472 => X"00000000",
    3473 => X"0000d1b7",
    3474 => X"00000256",
    3475 => X"000000fa",
    3476 => X"00000000",
    3477 => X"0000d1b7",
    3478 => X"0000024e",
    3479 => X"000000fa",
    3480 => X"00000000",
    3481 => X"0000d1b7",
    3482 => X"00000245",
    3483 => X"000000fa",
    3484 => X"00000000",
    3485 => X"0000d1b7",
    3486 => X"0000023d",
    3487 => X"000000fa",
    3488 => X"00000000",
    3489 => X"0000d1b7",
    3490 => X"00000235",
    3491 => X"000000fa",
    3492 => X"00000000",
    3493 => X"0000d1b7",
    3494 => X"0000022c",
    3495 => X"000000fa",
    3496 => X"00000000",
    3497 => X"0000d1b7",
    3498 => X"00000224",
    3499 => X"000000fa",
    3500 => X"00000000",
    3501 => X"0000d1b7",
    3502 => X"0000021c",
    3503 => X"000000fa",
    3504 => X"00000000",
    3505 => X"0000d1b7",
    3506 => X"00000214",
    3507 => X"000000fa",
    3508 => X"00000000",
    3509 => X"0000d1b7",
    3510 => X"0000020b",
    3511 => X"000000fa",
    3512 => X"00000000",
    3513 => X"0000d1b7",
    3514 => X"00000203",
    3515 => X"000000fa",
    3516 => X"00000000",
    3517 => X"0000d1b7",
    3518 => X"000001fb",
    3519 => X"000000fa",
    3520 => X"00000000",
    3521 => X"0000d1b7",
    3522 => X"000001f3",
    3523 => X"000000fa",
    3524 => X"00000000",
    3525 => X"0000d1b7",
    3526 => X"000001ec",
    3527 => X"000000fa",
    3528 => X"00000000",
    3529 => X"0000d1b7",
    3530 => X"000001e4",
    3531 => X"000000fa",
    3532 => X"00000000",
    3533 => X"0000d1b7",
    3534 => X"000001dc",
    3535 => X"000000fa",
    3536 => X"00000000",
    3537 => X"0000d1b7",
    3538 => X"000001d4",
    3539 => X"000000fa",
    3540 => X"00000000",
    3541 => X"0000d1b7",
    3542 => X"000001cc",
    3543 => X"000000fa",
    3544 => X"00000000",
    3545 => X"0000d1b7",
    3546 => X"000001c5",
    3547 => X"000000fa",
    3548 => X"00000000",
    3549 => X"0000d1b7",
    3550 => X"000001bd",
    3551 => X"000000fa",
    3552 => X"00000000",
    3553 => X"0000d1b7",
    3554 => X"000001b6",
    3555 => X"000000fa",
    3556 => X"00000000",
    3557 => X"0000d1b7",
    3558 => X"000001ae",
    3559 => X"000000fa",
    3560 => X"00000000",
    3561 => X"0000d1b7",
    3562 => X"000001a7",
    3563 => X"000000fa",
    3564 => X"00000000",
    3565 => X"0000d1b7",
    3566 => X"000001a0",
    3567 => X"000000fa",
    3568 => X"00000000",
    3569 => X"0000d1b7",
    3570 => X"00000198",
    3571 => X"000000fa",
    3572 => X"00000000",
    3573 => X"0000d1b7",
    3574 => X"00000191",
    3575 => X"000000fa",
    3576 => X"00000000",
    3577 => X"0000d1b7",
    3578 => X"0000018a",
    3579 => X"000000fa",
    3580 => X"00000000",
    3581 => X"0000d1b7",
    3582 => X"00000183",
    3583 => X"000000fa",
    3584 => X"00000000",
    3585 => X"0000d1b7",
    3586 => X"0000017c",
    3587 => X"000000fa",
    3588 => X"00000000",
    3589 => X"0000d1b7",
    3590 => X"00000175",
    3591 => X"000000fa",
    3592 => X"00000000",
    3593 => X"0000d1b7",
    3594 => X"0000016e",
    3595 => X"000000fa",
    3596 => X"00000000",
    3597 => X"0000d1b7",
    3598 => X"00000167",
    3599 => X"000000fa",
    3600 => X"00000000",
    3601 => X"0000d1b7",
    3602 => X"00000160",
    3603 => X"000000fa",
    3604 => X"00000000",
    3605 => X"0000d1b7",
    3606 => X"00000159",
    3607 => X"000000fa",
    3608 => X"00000000",
    3609 => X"0000d1b7",
    3610 => X"00000152",
    3611 => X"000000fa",
    3612 => X"00000000",
    3613 => X"0000d1b7",
    3614 => X"0000014c",
    3615 => X"000000fa",
    3616 => X"00000000",
    3617 => X"0000d1b7",
    3618 => X"00000145",
    3619 => X"000000fa",
    3620 => X"00000000",
    3621 => X"0000d1b7",
    3622 => X"0000013f",
    3623 => X"000000fa",
    3624 => X"00000000",
    3625 => X"0000d1b7",
    3626 => X"00000138",
    3627 => X"000000fa",
    3628 => X"00000000",
    3629 => X"0000d1b7",
    3630 => X"00000132",
    3631 => X"000000fa",
    3632 => X"00000000",
    3633 => X"0000d1b7",
    3634 => X"0000012b",
    3635 => X"000000fa",
    3636 => X"00000000",
    3637 => X"0000d1b7",
    3638 => X"00000125",
    3639 => X"000000fa",
    3640 => X"00000000",
    3641 => X"0000d1b7",
    3642 => X"0000011f",
    3643 => X"000000fa",
    3644 => X"00000000",
    3645 => X"0000d1b7",
    3646 => X"00000119",
    3647 => X"000000fa",
    3648 => X"00000000",
    3649 => X"0000d1b7",
    3650 => X"00000113",
    3651 => X"000000fa",
    3652 => X"00000000",
    3653 => X"0000d1b7",
    3654 => X"0000010d",
    3655 => X"000000fa",
    3656 => X"00000000",
    3657 => X"0000d1b7",
    3658 => X"00000107",
    3659 => X"000000fa",
    3660 => X"00000000",
    3661 => X"0000d1b7",
    3662 => X"00000101",
    3663 => X"000000fa",
    3664 => X"00000000",
    3665 => X"0000d1b7",
    3666 => X"000000fb",
    3667 => X"000000fa",
    3668 => X"00000000",
    3669 => X"0000d1b7",
    3670 => X"000000f5",
    3671 => X"000000fa",
    3672 => X"00000000",
    3673 => X"0000d1b7",
    3674 => X"000000ef",
    3675 => X"000000fa",
    3676 => X"00000000",
    3677 => X"0000d1b7",
    3678 => X"000000ea",
    3679 => X"000000fa",
    3680 => X"00000000",
    3681 => X"0000d1b7",
    3682 => X"000000e4",
    3683 => X"000000fa",
    3684 => X"00000000",
    3685 => X"0000d1b7",
    3686 => X"000000de",
    3687 => X"000000fa",
    3688 => X"00000000",
    3689 => X"0000d1b7",
    3690 => X"000000d9",
    3691 => X"000000fa",
    3692 => X"00000000",
    3693 => X"0000d1b7",
    3694 => X"000000d3",
    3695 => X"000000fa",
    3696 => X"00000000",
    3697 => X"0000d1b7",
    3698 => X"000000ce",
    3699 => X"000000fa",
    3700 => X"00000000",
    3701 => X"0000d1b7",
    3702 => X"000000c9",
    3703 => X"000000fa",
    3704 => X"00000000",
    3705 => X"0000d1b7",
    3706 => X"000000c4",
    3707 => X"000000fa",
    3708 => X"00000000",
    3709 => X"0000d1b7",
    3710 => X"000000be",
    3711 => X"000000fa",
    3712 => X"00000000",
    3713 => X"0000d1b7",
    3714 => X"000000b9",
    3715 => X"000000fa",
    3716 => X"00000000",
    3717 => X"0000d1b7",
    3718 => X"000000b4",
    3719 => X"000000fa",
    3720 => X"00000000",
    3721 => X"0000d1b7",
    3722 => X"000000af",
    3723 => X"000000fa",
    3724 => X"00000000",
    3725 => X"0000d1b7",
    3726 => X"000000aa",
    3727 => X"000000fa",
    3728 => X"00000000",
    3729 => X"0000d1b7",
    3730 => X"000000a6",
    3731 => X"000000fa",
    3732 => X"00000000",
    3733 => X"0000d1b7",
    3734 => X"000000a1",
    3735 => X"000000fa",
    3736 => X"00000000",
    3737 => X"0000d1b7",
    3738 => X"0000009c",
    3739 => X"000000fa",
    3740 => X"00000000",
    3741 => X"0000d1b7",
    3742 => X"00000098",
    3743 => X"000000fa",
    3744 => X"00000000",
    3745 => X"0000d1b7",
    3746 => X"00000093",
    3747 => X"000000fa",
    3748 => X"00000000",
    3749 => X"0000d1b7",
    3750 => X"0000008e",
    3751 => X"000000fa",
    3752 => X"00000000",
    3753 => X"0000d1b7",
    3754 => X"0000008a",
    3755 => X"000000fa",
    3756 => X"00000000",
    3757 => X"0000d1b7",
    3758 => X"00000086",
    3759 => X"000000fa",
    3760 => X"00000000",
    3761 => X"0000d1b7",
    3762 => X"00000081",
    3763 => X"000000fa",
    3764 => X"00000000",
    3765 => X"0000d1b7",
    3766 => X"0000007d",
    3767 => X"000000fa",
    3768 => X"00000000",
    3769 => X"0000d1b7",
    3770 => X"00000079",
    3771 => X"000000fa",
    3772 => X"00000000",
    3773 => X"0000d1b7",
    3774 => X"00000075",
    3775 => X"000000fa",
    3776 => X"00000000",
    3777 => X"0000d1b7",
    3778 => X"00000071",
    3779 => X"000000fa",
    3780 => X"00000000",
    3781 => X"0000d1b7",
    3782 => X"0000006d",
    3783 => X"000000fa",
    3784 => X"00000000",
    3785 => X"0000d1b7",
    3786 => X"00000069",
    3787 => X"000000fa",
    3788 => X"00000000",
    3789 => X"0000d1b7",
    3790 => X"00000065",
    3791 => X"000000fa",
    3792 => X"00000000",
    3793 => X"0000d1b7",
    3794 => X"00000061",
    3795 => X"000000fa",
    3796 => X"00000000",
    3797 => X"0000d1b7",
    3798 => X"0000005e",
    3799 => X"000000fa",
    3800 => X"00000000",
    3801 => X"0000d1b7",
    3802 => X"0000005a",
    3803 => X"000000fa",
    3804 => X"00000000",
    3805 => X"0000d1b7",
    3806 => X"00000057",
    3807 => X"000000fa",
    3808 => X"00000000",
    3809 => X"0000d1b7",
    3810 => X"00000053",
    3811 => X"000000fa",
    3812 => X"00000000",
    3813 => X"0000d1b7",
    3814 => X"00000050",
    3815 => X"000000fa",
    3816 => X"00000000",
    3817 => X"0000d1b7",
    3818 => X"0000004c",
    3819 => X"000000fa",
    3820 => X"00000000",
    3821 => X"0000d1b7",
    3822 => X"00000049",
    3823 => X"000000fa",
    3824 => X"00000000",
    3825 => X"0000d1b7",
    3826 => X"00000046",
    3827 => X"000000fa",
    3828 => X"00000000",
    3829 => X"0000d1b7",
    3830 => X"00000043",
    3831 => X"000000fa",
    3832 => X"00000000",
    3833 => X"0000d1b7",
    3834 => X"00000040",
    3835 => X"000000fa",
    3836 => X"00000000",
    3837 => X"0000d1b7",
    3838 => X"0000003d",
    3839 => X"000000fa",
    3840 => X"00000000",
    3841 => X"0000d1b7",
    3842 => X"0000003a",
    3843 => X"000000fa",
    3844 => X"00000000",
    3845 => X"0000d1b7",
    3846 => X"00000037",
    3847 => X"000000fa",
    3848 => X"00000000",
    3849 => X"0000d1b7",
    3850 => X"00000034",
    3851 => X"000000fa",
    3852 => X"00000000",
    3853 => X"0000d1b7",
    3854 => X"00000032",
    3855 => X"000000fa",
    3856 => X"00000000",
    3857 => X"0000d1b7",
    3858 => X"0000002f",
    3859 => X"000000fa",
    3860 => X"00000000",
    3861 => X"0000d1b7",
    3862 => X"0000002c",
    3863 => X"000000fa",
    3864 => X"00000000",
    3865 => X"0000d1b7",
    3866 => X"0000002a",
    3867 => X"000000fa",
    3868 => X"00000000",
    3869 => X"0000d1b7",
    3870 => X"00000027",
    3871 => X"000000fa",
    3872 => X"00000000",
    3873 => X"0000d1b7",
    3874 => X"00000025",
    3875 => X"000000fa",
    3876 => X"00000000",
    3877 => X"0000d1b7",
    3878 => X"00000023",
    3879 => X"000000fa",
    3880 => X"00000000",
    3881 => X"0000d1b7",
    3882 => X"00000021",
    3883 => X"000000fa",
    3884 => X"00000000",
    3885 => X"0000d1b7",
    3886 => X"0000001f",
    3887 => X"000000fa",
    3888 => X"00000000",
    3889 => X"0000d1b7",
    3890 => X"0000001c",
    3891 => X"000000fa",
    3892 => X"00000000",
    3893 => X"0000d1b7",
    3894 => X"0000001a",
    3895 => X"000000fa",
    3896 => X"00000000",
    3897 => X"0000d1b7",
    3898 => X"00000019",
    3899 => X"000000fa",
    3900 => X"00000000",
    3901 => X"0000d1b7",
    3902 => X"00000017",
    3903 => X"000000fa",
    3904 => X"00000000",
    3905 => X"0000d1b7",
    3906 => X"00000015",
    3907 => X"000000fa",
    3908 => X"00000000",
    3909 => X"0000d1b7",
    3910 => X"00000013",
    3911 => X"000000fa",
    3912 => X"00000000",
    3913 => X"0000d1b7",
    3914 => X"00000012",
    3915 => X"000000fa",
    3916 => X"00000000",
    3917 => X"0000d1b7",
    3918 => X"00000010",
    3919 => X"000000fa",
    3920 => X"00000000",
    3921 => X"0000d1b7",
    3922 => X"0000000f",
    3923 => X"000000fa",
    3924 => X"00000000",
    3925 => X"0000d1b7",
    3926 => X"0000000d",
    3927 => X"000000fa",
    3928 => X"00000000",
    3929 => X"0000d1b7",
    3930 => X"0000000c",
    3931 => X"000000fa",
    3932 => X"00000000",
    3933 => X"0000d1b7",
    3934 => X"0000000b",
    3935 => X"000000fa",
    3936 => X"00000000",
    3937 => X"0000d1b7",
    3938 => X"00000009",
    3939 => X"000000fa",
    3940 => X"00000000",
    3941 => X"0000d1b7",
    3942 => X"00000008",
    3943 => X"000000fa",
    3944 => X"00000000",
    3945 => X"0000d1b7",
    3946 => X"00000007",
    3947 => X"000000fa",
    3948 => X"00000000",
    3949 => X"0000d1b7",
    3950 => X"00000006",
    3951 => X"000000fa",
    3952 => X"00000000",
    3953 => X"0000d1b7",
    3954 => X"00000005",
    3955 => X"000000fa",
    3956 => X"00000000",
    3957 => X"0000d1b7",
    3958 => X"00000004",
    3959 => X"000000fa",
    3960 => X"00000000",
    3961 => X"0000d1b7",
    3962 => X"00000004",
    3963 => X"000000fa",
    3964 => X"00000000",
    3965 => X"0000d1b7",
    3966 => X"00000003",
    3967 => X"000000fa",
    3968 => X"00000000",
    3969 => X"0000d1b7",
    3970 => X"00000002",
    3971 => X"000000fa",
    3972 => X"00000000",
    3973 => X"0000d1b7",
    3974 => X"00000002",
    3975 => X"000000fa",
    3976 => X"00000000",
    3977 => X"0000d1b7",
    3978 => X"00000001",
    3979 => X"000000fa",
    3980 => X"00000000",
    3981 => X"0000d1b7",
    3982 => X"00000001",
    3983 => X"000000fa",
    3984 => X"00000000",
    3985 => X"0000d1b7",
    3986 => X"00000001",
    3987 => X"000000fa",
    3988 => X"00000000",
    3989 => X"0000d1b7",
    3990 => X"00000000",
    3991 => X"000000fa",
    3992 => X"00000000",
    3993 => X"0000d1b7",
    3994 => X"00000000",
    3995 => X"000000fa",
    3996 => X"00000000",
    3997 => X"0000d1b7",
    3998 => X"00000000",
    3999 => X"000000fa",
    4000 => X"00000000",
    4001 => X"0000d1b7",
    4002 => X"00000000",
    4003 => X"000003e8",
    4004 => X"00000000",
    4005 => X"0000d1b7",
    4006 => X"00000000",
    4007 => X"00000000");
end DataPackage;
